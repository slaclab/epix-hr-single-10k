------------------------------------------------------------------------------
-- This file is part of 'EPIX Development Firmware'.
-- It is subject to the license terms in the LICENSE.txt file found in the 
-- top-level directory of this distribution and at: 
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html. 
-- No part of 'EPIX Development Firmware', including this file, 
-- may be copied, modified, propagated, or distributed except according to 
-- the terms contained in the LICENSE.txt file.
------------------------------------------------------------------------------
-- Auto-generated package containing LUT initialization data
-- for conversion of the environmental data of the EPIX detector
-- To regenerate use envDataFpgaLut.cpp
-- Maciej Kwiatkowski (mkwiatko@slac.stanford.edu)
-- Generation date 12/03/2015

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

package SlowAdcPkg is
constant INIT_H_TH0_00 : bit_vector(255 downto 0) := X"2626262626262626262626262626262626262626262626262626262626262626";
constant INIT_L_TH0_00 : bit_vector(255 downto 0) := X"016FE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1";
constant INIT_H_TH0_01 : bit_vector(255 downto 0) := X"1D1D1D1D1E1E1E1E1E1F1F1F1F20202020212121212222222323232424242525";
constant INIT_L_TH0_01 : bit_vector(255 downto 0) := X"4070A1D306396EA4DB134C87C3003F7FC1044A90D92471C01165BB1470D03298";
constant INIT_H_TH0_02 : bit_vector(255 downto 0) := X"1818181819191919191919191A1A1A1A1A1A1A1B1B1B1B1B1B1C1C1C1C1C1C1D";
constant INIT_L_TH0_02 : bit_vector(255 downto 0) := X"98B6D4F21131507091B2D3F5183B5E82A6CBF1173D648CB5DE07325D89B5E311";
constant INIT_H_TH0_03 : bit_vector(255 downto 0) := X"1515151515151516161616161616161616161717171717171717171818181818";
constant INIT_L_TH0_03 : bit_vector(255 downto 0) := X"788DA3B8CEE4FB11283F566E859DB5CEE7FF19324C66809BB5D1EC0824405D7A";
constant INIT_H_TH0_04 : bit_vector(255 downto 0) := X"1313131313131313131313131314141414141414141414141414141515151515";
constant INIT_L_TH0_04 : bit_vector(255 downto 0) := X"2334445566778899ABBCCEDFF10316283A4D60738699ACC0D4E8FC1024394E63";
constant INIT_H_TH0_05 : bit_vector(255 downto 0) := X"1111111111111111111111111111121212121212121212121212121212121313";
constant INIT_L_TH0_05 : bit_vector(255 downto 0) := X"4B586673818E9CAAB8C6D4E2F1FF0D1C2B39485766758594A4B3C3D3E3F30313";
constant INIT_H_TH0_06 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F1010101010101010101010101010101010101010101111111111";
constant INIT_L_TH0_06 : bit_vector(255 downto 0) := X"C5D0DCE7F2FE0915202C38434F5B67737F8C98A4B0BDC9D6E3EFFC091623303E";
constant INIT_H_TH0_07 : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_TH0_07 : bit_vector(255 downto 0) := X"7B848E98A1ABB5BFC9D3DDE7F1FB050F1A242E39434E58636E78838E99A4AFBA";
constant INIT_H_TH0_08 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_TH0_08 : bit_vector(255 downto 0) := X"5C656D767E878F98A0A9B2BAC3CCD5DEE7F0F9020B141D262F39424B555E6871";
constant INIT_H_TH0_09 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_TH0_09 : bit_vector(255 downto 0) := X"60686F777E868D959DA4ACB4BBC3CBD3DBE2EAF2FA020A121A232B333B434C54";
constant INIT_H_TH0_0A : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_TH0_0A : bit_vector(255 downto 0) := X"80868D949AA1A8AFB6BCC3CAD1D8DFE6EDF4FB020910171F262D343C434A5259";
constant INIT_H_TH0_0B : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_TH0_0B : bit_vector(255 downto 0) := X"B5BBC1C7CDD3DAE0E6ECF2F8FF050B11181E242B31383E454B52585F656C7279";
constant INIT_H_TH0_0C : bit_vector(255 downto 0) := X"090A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_TH0_0C : bit_vector(255 downto 0) := X"FD02080D13191E24292F353A40464B51575D62686E747A7F858B91979DA3A9AF";
constant INIT_H_TH0_0D : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_TH0_0D : bit_vector(255 downto 0) := X"54595E63686E73787D82878C92979CA1A7ACB1B7BCC1C7CCD1D7DCE1E7ECF2F7";
constant INIT_H_TH0_0E : bit_vector(255 downto 0) := X"0808080808080808080808080808080909090909090909090909090909090909";
constant INIT_L_TH0_0E : bit_vector(255 downto 0) := X"B9BDC2C7CBD0D5DADEE3E8EDF1F6FB00050A0F13181D22272C31363B40454A4F";
constant INIT_H_TH0_0F : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_TH0_0F : bit_vector(255 downto 0) := X"282D31353A3E43474B5054595D62666B6F74787D81868A8F93989DA1A6ABAFB4";
constant INIT_H_TH0_10 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707080808080808080808";
constant INIT_L_TH0_10 : bit_vector(255 downto 0) := X"A2A6AAAEB2B6BBBFC3C7CBCFD3D7DCE0E4E8ECF1F5F9FD02060A0E13171B2024";
constant INIT_H_TH0_11 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_TH0_11 : bit_vector(255 downto 0) := X"24282C3034383B3F43474B4F53565A5E62666A6E72767A7E82868A8E92969A9E";
constant INIT_H_TH0_12 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606070707070707070707";
constant INIT_L_TH0_12 : bit_vector(255 downto 0) := X"AEB2B6B9BDC0C4C8CBCFD3D6DADEE1E5E9ECF0F4F7FBFF03060A0E1215191D21";
constant INIT_H_TH0_13 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_TH0_13 : bit_vector(255 downto 0) := X"3F43464A4D5054575B5E6165686C6F73767A7D8184888B8F9296999DA0A4A7AB";
constant INIT_H_TH0_14 : bit_vector(255 downto 0) := X"0505050505050505050505050506060606060606060606060606060606060606";
constant INIT_L_TH0_14 : bit_vector(255 downto 0) := X"D6DADDE0E3E6EAEDF0F3F7FAFD0004070A0D1114171B1E2125282B2F3235393C";
constant INIT_H_TH0_15 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_TH0_15 : bit_vector(255 downto 0) := X"7376797C7F8285888B8E9195989B9EA1A4A7AAADB0B4B7BABDC0C3C6CACDD0D3";
constant INIT_H_TH0_16 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_TH0_16 : bit_vector(255 downto 0) := X"14171A1D202326292C2F3134373A3D404346494C4F5255585B5E6164676A6D70";
constant INIT_H_TH0_17 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040405050505050505";
constant INIT_L_TH0_17 : bit_vector(255 downto 0) := X"BBBDC0C3C6C8CBCED1D3D6D9DCDFE1E4E7EAEDEFF2F5F8FBFE000306090C0F12";
constant INIT_H_TH0_18 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_TH0_18 : bit_vector(255 downto 0) := X"65676A6D6F7275777A7C7F8284878A8C8F9295979A9D9FA2A5A7AAADB0B2B5B8";
constant INIT_H_TH0_19 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_TH0_19 : bit_vector(255 downto 0) := X"1315181A1D1F222427292C2F313436393B3E404346484B4D505255585A5D5F62";
constant INIT_H_TH0_1A : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030304040404040404";
constant INIT_L_TH0_1A : bit_vector(255 downto 0) := X"C4C7C9CBCED0D3D5D8DADCDFE1E4E6E9EBEEF0F2F5F7FAFCFF010406090B0E10";
constant INIT_H_TH0_1B : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_TH0_1B : bit_vector(255 downto 0) := X"797B7E80828587898B8E909295979A9C9EA1A3A5A8AAACAFB1B3B6B8BBBDBFC2";
constant INIT_H_TH0_1C : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_TH0_1C : bit_vector(255 downto 0) := X"313335373A3C3E40424547494B4E50525457595B5D60626467696B6D70727477";
constant INIT_H_TH0_1D : bit_vector(255 downto 0) := X"0202020202020202020203030303030303030303030303030303030303030303";
constant INIT_L_TH0_1D : bit_vector(255 downto 0) := X"EBEDEFF2F4F6F8FAFCFE01030507090B0E10121416181B1D1F212326282A2C2E";
constant INIT_H_TH0_1E : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_TH0_1E : bit_vector(255 downto 0) := X"A8AAACAEB0B2B4B7B9BBBDBFC1C3C5C7C9CBCDD0D2D4D6D8DADCDEE0E3E5E7E9";
constant INIT_H_TH0_1F : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_TH0_1F : bit_vector(255 downto 0) := X"686A6C6D6F71737577797B7D7F818486888A8C8E90929496989A9C9EA0A2A4A6";
constant INIT_H_TH0_20 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_TH0_20 : bit_vector(255 downto 0) := X"292B2D2F31333537393B3C3E40424446484A4C4E50525456585A5C5E60626466";
constant INIT_H_TH0_21 : bit_vector(255 downto 0) := X"0101010101010101010102020202020202020202020202020202020202020202";
constant INIT_L_TH0_21 : bit_vector(255 downto 0) := X"EDEFF1F3F4F6F8FAFCFE0001030507090B0D0F10121416181A1C1E2022232527";
constant INIT_H_TH0_22 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_TH0_22 : bit_vector(255 downto 0) := X"B3B4B6B8BABCBDBFC1C3C5C6C8CACCCED0D1D3D5D7D9DBDCDEE0E2E4E6E7E9EB";
constant INIT_H_TH0_23 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_TH0_23 : bit_vector(255 downto 0) := X"7A7C7E7F81838586888A8C8D8F91939496989A9C9D9FA1A3A4A6A8AAACADAFB1";
constant INIT_H_TH0_24 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_TH0_24 : bit_vector(255 downto 0) := X"444547494A4C4E4F51535456585A5B5D5F6062646667696B6C6E707273757778";
constant INIT_H_TH0_25 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_TH0_25 : bit_vector(255 downto 0) := X"0E1012131517181A1C1D1F2122242527292A2C2E2F3133343638393B3D3E4042";
constant INIT_H_TH0_26 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000010101010101010101";
constant INIT_L_TH0_26 : bit_vector(255 downto 0) := X"DBDDDEE0E1E3E5E6E8E9EBEDEEF0F1F3F5F6F8F9FBFDFE0001030506080A0B0D";
constant INIT_H_TH0_27 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_TH0_27 : bit_vector(255 downto 0) := X"A9AAACAEAFB1B2B4B5B7B8BABCBDBFC0C2C3C5C6C8CACBCDCED0D1D3D5D6D8D9";
constant INIT_H_TH0_28 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_TH0_28 : bit_vector(255 downto 0) := X"787A7B7D7E808183848687898A8C8D8F9092939597989A9B9D9EA0A1A3A4A6A7";
constant INIT_H_TH0_29 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_TH0_29 : bit_vector(255 downto 0) := X"494A4C4D4F505253555658595B5C5E5F606263656668696B6C6E6F7172747577";
constant INIT_H_TH0_2A : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_TH0_2A : bit_vector(255 downto 0) := X"1B1C1E1F212223252628292B2C2D2F303233353638393A3C3D3F404243454648";
constant INIT_H_TH0_2B : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000";
constant INIT_L_TH0_2B : bit_vector(255 downto 0) := X"EEEFF1F2F4F5F6F8F9FBFCFDFF000103040607090A0B0D0E1011121415171819";
constant INIT_H_TH0_2C : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_TH0_2C : bit_vector(255 downto 0) := X"C2C4C5C6C8C9CACCCDCED0D1D3D4D5D7D8D9DBDCDDDFE0E2E3E4E6E7E8EAEBED";
constant INIT_H_TH0_2D : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_TH0_2D : bit_vector(255 downto 0) := X"98999A9C9D9E9FA1A2A3A5A6A7A9AAABADAEAFB1B2B3B5B6B7B9BABCBDBEC0C1";
constant INIT_H_TH0_2E : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_TH0_2E : bit_vector(255 downto 0) := X"6E6F707273747677787A7B7C7D7F80818384858788898A8C8D8E909192949596";
constant INIT_H_TH0_2F : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_TH0_2F : bit_vector(255 downto 0) := X"454748494A4C4D4E4F51525354565758595B5C5D5F60616264656668696A6B6D";
constant INIT_H_TH0_30 : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_TH0_30 : bit_vector(255 downto 0) := X"1E1F20212224252627292A2B2C2E2F30313334353638393A3B3C3E3F40424344";
constant INIT_H_TH0_31 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_TH0_31 : bit_vector(255 downto 0) := X"F7F8F9FAFCFDFEFF00020304050608090A0B0C0E0F10111314151617191A1B1C";
constant INIT_H_TH0_32 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH0_32 : bit_vector(255 downto 0) := X"D1D2D3D4D5D7D8D9DADBDDDEDFE0E1E2E4E5E6E7E8EAEBECEDEEF0F1F2F3F4F6";
constant INIT_H_TH0_33 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH0_33 : bit_vector(255 downto 0) := X"ACADAEAFB0B1B3B4B5B6B7B8B9BBBCBDBEBFC0C2C3C4C5C6C7C9CACBCCCDCED0";
constant INIT_H_TH0_34 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH0_34 : bit_vector(255 downto 0) := X"87888A8B8C8D8E8F9091939495969798999B9C9D9E9FA0A1A2A4A5A6A7A8A9AB";
constant INIT_H_TH0_35 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH0_35 : bit_vector(255 downto 0) := X"6465666768696A6B6D6E6F7071727374757778797A7B7C7D7E7F818283848586";
constant INIT_H_TH0_36 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH0_36 : bit_vector(255 downto 0) := X"41424344454647484A4B4C4D4E4F5051525354565758595A5B5C5D5E5F606263";
constant INIT_H_TH0_37 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH0_37 : bit_vector(255 downto 0) := X"1F202122232425262728292A2B2D2E2F303132333435363738393A3C3D3E3F40";
constant INIT_H_TH0_38 : bit_vector(255 downto 0) := X"FDFDFDFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH0_38 : bit_vector(255 downto 0) := X"FDFEFF0001030405060708090A0B0C0D0E0F1011121314151617181A1B1C1D1E";
constant INIT_H_TH0_39 : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH0_39 : bit_vector(255 downto 0) := X"DDDEDFE0E1E2E3E4E5E6E7E8E9EAEBECEDEEEFF0F1F2F3F4F5F6F7F8F9FAFBFC";
constant INIT_H_TH0_3A : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH0_3A : bit_vector(255 downto 0) := X"BCBDBEBFC0C1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADB";
constant INIT_H_TH0_3B : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH0_3B : bit_vector(255 downto 0) := X"9D9E9FA0A1A2A3A4A5A6A7A8A9AAABABACADAEAFB0B1B2B3B4B5B6B7B8B9BABB";
constant INIT_H_TH0_3C : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH0_3C : bit_vector(255 downto 0) := X"7E7F80818283848585868788898A8B8C8D8E8F909192939495969798999A9B9C";
constant INIT_H_TH0_3D : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH0_3D : bit_vector(255 downto 0) := X"5F606162636465666768696A6B6C6D6E6F6F707172737475767778797A7B7C7D";
constant INIT_H_TH0_3E : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH0_3E : bit_vector(255 downto 0) := X"4142434445464748494A4B4C4D4E4E4F505152535455565758595A5B5C5D5D5E";
constant INIT_H_TH0_3F : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH0_3F : bit_vector(255 downto 0) := X"2425262728292A2B2B2C2D2E2F30313233343536363738393A3B3C3D3E3F4041";
constant INIT_H_TH0_40 : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH0_40 : bit_vector(255 downto 0) := X"0708090A0B0C0D0E0E0F10111213141516171718191A1B1C1D1E1F2021212223";
constant INIT_H_TH0_41 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFDFDFDFDFDFDFDFD";
constant INIT_L_TH0_41 : bit_vector(255 downto 0) := X"EBECEDEEEEEFF0F1F2F3F4F5F6F6F7F8F9FAFBFCFDFEFEFF0001020304050606";
constant INIT_H_TH0_42 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH0_42 : bit_vector(255 downto 0) := X"CFD0D1D2D3D3D4D5D6D7D8D9D9DADBDCDDDEDFE0E0E1E2E3E4E5E6E7E7E8E9EA";
constant INIT_H_TH0_43 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH0_43 : bit_vector(255 downto 0) := X"B4B5B5B6B7B8B9BABBBBBCBDBEBFC0C0C1C2C3C4C5C6C6C7C8C9CACBCCCDCDCE";
constant INIT_H_TH0_44 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH0_44 : bit_vector(255 downto 0) := X"999A9A9B9C9D9E9F9FA0A1A2A3A4A4A5A6A7A8A9AAAAABACADAEAFAFB0B1B2B3";
constant INIT_H_TH0_45 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH0_45 : bit_vector(255 downto 0) := X"7E7F8081828283848586868788898A8B8B8C8D8E8F9090919293949595969798";
constant INIT_H_TH0_46 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH0_46 : bit_vector(255 downto 0) := X"646566676768696A6B6B6C6D6E6F6F7071727374747576777878797A7B7C7D7D";
constant INIT_H_TH0_47 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH0_47 : bit_vector(255 downto 0) := X"4A4B4C4D4E4E4F5051525253545556565758595A5A5B5C5D5E5E5F6061626363";
constant INIT_H_TH0_48 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH0_48 : bit_vector(255 downto 0) := X"31323333343536373738393A3B3B3C3D3E3F3F4041424243444546464748494A";
constant INIT_H_TH0_49 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH0_49 : bit_vector(255 downto 0) := X"18191A1B1B1C1D1E1E1F202122222324252526272829292A2B2C2C2D2E2F3030";
constant INIT_H_TH0_4A : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH0_4A : bit_vector(255 downto 0) := X"000001020303040506070708090A0A0B0C0D0D0E0F1011111213141415161717";
constant INIT_H_TH0_4B : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH0_4B : bit_vector(255 downto 0) := X"E8E8E9EAEBEBECEDEEEEEFF0F1F1F2F3F4F4F5F6F7F7F8F9FAFAFBFCFDFDFEFF";
constant INIT_H_TH0_4C : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH0_4C : bit_vector(255 downto 0) := X"D0D0D1D2D3D3D4D5D6D6D7D8D9D9DADBDCDCDDDEDFDFE0E1E2E2E3E4E5E5E6E7";
constant INIT_H_TH0_4D : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH0_4D : bit_vector(255 downto 0) := X"B8B9BABABBBCBDBDBEBFC0C0C1C2C2C3C4C5C5C6C7C8C8C9CACBCBCCCDCDCECF";
constant INIT_H_TH0_4E : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH0_4E : bit_vector(255 downto 0) := X"A1A2A3A3A4A5A5A6A7A8A8A9AAAAABACADADAEAFB0B0B1B2B2B3B4B5B5B6B7B7";
constant INIT_H_TH0_4F : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH0_4F : bit_vector(255 downto 0) := X"8A8B8C8C8D8E8F8F90919192939494959696979898999A9B9B9C9D9E9E9FA0A0";
constant INIT_H_TH0_50 : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH0_50 : bit_vector(255 downto 0) := X"7474757677777879797A7B7B7C7D7E7E7F80808182838384858586878788898A";
constant INIT_H_TH0_51 : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH0_51 : bit_vector(255 downto 0) := X"5E5E5F6060616262636464656667676869696A6B6B6C6D6E6E6F707071727273";
constant INIT_H_TH0_52 : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH0_52 : bit_vector(255 downto 0) := X"4848494A4A4B4C4C4D4E4F4F5051515253535455555657575859595A5B5C5C5D";
constant INIT_H_TH0_53 : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH0_53 : bit_vector(255 downto 0) := X"32333334353536373738393A3A3B3C3C3D3E3E3F404041424243444445464647";
constant INIT_H_TH0_54 : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH0_54 : bit_vector(255 downto 0) := X"1D1D1E1F1F2021212223232425252627272829292A2B2B2C2D2D2E2F2F303131";
constant INIT_H_TH0_55 : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH0_55 : bit_vector(255 downto 0) := X"0808090A0A0B0C0C0D0E0E0F1010111212131414151616171818191A1A1B1B1C";
constant INIT_H_TH0_56 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH0_56 : bit_vector(255 downto 0) := X"F3F4F4F5F6F6F7F8F8F9F9FAFBFBFCFDFDFEFFFF000101020303040505060607";
constant INIT_H_TH0_57 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_57 : bit_vector(255 downto 0) := X"DFDFE0E0E1E2E2E3E4E4E5E6E6E7E7E8E9E9EAEBEBECEDEDEEEFEFF0F0F1F2F2";
constant INIT_H_TH0_58 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_58 : bit_vector(255 downto 0) := X"CACBCCCCCDCDCECFCFD0D1D1D2D2D3D4D4D5D6D6D7D8D8D9D9DADBDBDCDDDDDE";
constant INIT_H_TH0_59 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_59 : bit_vector(255 downto 0) := X"B6B7B8B8B9B9BABBBBBCBDBDBEBEBFC0C0C1C2C2C3C3C4C5C5C6C7C7C8C8C9CA";
constant INIT_H_TH0_5A : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_5A : bit_vector(255 downto 0) := X"A3A3A4A4A5A6A6A7A7A8A9A9AAABABACACADAEAEAFB0B0B1B1B2B3B3B4B4B5B6";
constant INIT_H_TH0_5B : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_5B : bit_vector(255 downto 0) := X"8F90909192929393949595969697989899999A9B9B9C9C9D9E9E9FA0A0A1A1A2";
constant INIT_H_TH0_5C : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_5C : bit_vector(255 downto 0) := X"7C7C7D7E7E7F7F808181828283848485858687878888898A8A8B8B8C8D8D8E8E";
constant INIT_H_TH0_5D : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_5D : bit_vector(255 downto 0) := X"69696A6B6B6C6C6D6E6E6F6F70717172727373747575767677787879797A7B7B";
constant INIT_H_TH0_5E : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_5E : bit_vector(255 downto 0) := X"5657575858595A5A5B5B5C5C5D5E5E5F5F606161626263636465656666676868";
constant INIT_H_TH0_5F : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_5F : bit_vector(255 downto 0) := X"43444545464647474849494A4A4B4C4C4D4D4E4E4F5050515152535354545555";
constant INIT_H_TH0_60 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_60 : bit_vector(255 downto 0) := X"3132323333343435363637373838393A3A3B3B3C3D3D3E3E3F3F404141424243";
constant INIT_H_TH0_61 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_61 : bit_vector(255 downto 0) := X"1F1F20212122222323242525262627272829292A2A2B2B2C2C2D2E2E2F2F3030";
constant INIT_H_TH0_62 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_62 : bit_vector(255 downto 0) := X"0D0E0E0F0F1010111112131314141515161617181819191A1A1B1C1C1D1D1E1E";
constant INIT_H_TH0_63 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH0_63 : bit_vector(255 downto 0) := X"FBFCFCFDFDFEFFFF0000010102020303040505060607070808090A0A0B0B0C0C";
constant INIT_H_TH0_64 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_64 : bit_vector(255 downto 0) := X"EAEAEBEBECECEDEDEEEFEFF0F0F1F1F2F2F3F3F4F5F5F6F6F7F7F8F8F9FAFAFB";
constant INIT_H_TH0_65 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_65 : bit_vector(255 downto 0) := X"D8D9D9DADADBDCDCDDDDDEDEDFDFE0E0E1E1E2E3E3E4E4E5E5E6E6E7E7E8E9E9";
constant INIT_H_TH0_66 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_66 : bit_vector(255 downto 0) := X"C7C8C8C9C9CACACBCBCCCCCDCECECFCFD0D0D1D1D2D2D3D3D4D5D5D6D6D7D7D8";
constant INIT_H_TH0_67 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_67 : bit_vector(255 downto 0) := X"B6B7B7B8B8B9B9BABABBBBBCBCBDBEBEBFBFC0C0C1C1C2C2C3C3C4C4C5C6C6C7";
constant INIT_H_TH0_68 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_68 : bit_vector(255 downto 0) := X"A5A6A6A7A7A8A8A9AAAAABABACACADADAEAEAFAFB0B0B1B1B2B2B3B3B4B5B5B6";
constant INIT_H_TH0_69 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_69 : bit_vector(255 downto 0) := X"959596969797989899999A9A9B9B9C9C9D9E9E9F9FA0A0A1A1A2A2A3A3A4A4A5";
constant INIT_H_TH0_6A : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_6A : bit_vector(255 downto 0) := X"84858586868787888889898A8A8B8B8C8C8D8D8E8F8F90909191929293939494";
constant INIT_H_TH0_6B : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_6B : bit_vector(255 downto 0) := X"74747575767777787879797A7A7B7B7C7C7D7D7E7E7F7F808081818282838384";
constant INIT_H_TH0_6C : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_6C : bit_vector(255 downto 0) := X"6464656566666767686869696A6A6B6B6C6C6D6D6E6E6F6F7070717172727373";
constant INIT_H_TH0_6D : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_6D : bit_vector(255 downto 0) := X"5454555556565757585859595A5A5B5B5C5C5D5D5E5E5F5F6060616162626363";
constant INIT_H_TH0_6E : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_6E : bit_vector(255 downto 0) := X"44454546464747484849494A4A4B4B4C4C4C4D4D4E4E4F4F5050515152525353";
constant INIT_H_TH0_6F : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_6F : bit_vector(255 downto 0) := X"35353536363737383839393A3A3B3B3C3C3D3D3E3E3F3F404041414242434344";
constant INIT_H_TH0_70 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_70 : bit_vector(255 downto 0) := X"252626262727282829292A2A2B2B2C2C2D2D2E2E2F2F30303131323233333434";
constant INIT_H_TH0_71 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_71 : bit_vector(255 downto 0) := X"16161717181819191A1A1A1B1B1C1C1D1D1E1E1F1F2020212122222323242425";
constant INIT_H_TH0_72 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_72 : bit_vector(255 downto 0) := X"070707080809090A0A0B0B0C0C0D0D0E0E0F0F10101011111212131314141515";
constant INIT_H_TH0_73 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH0_73 : bit_vector(255 downto 0) := X"F8F8F8F9F9FAFAFBFBFCFCFDFDFEFEFFFFFF0000010102020303040405050606";
constant INIT_H_TH0_74 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH0_74 : bit_vector(255 downto 0) := X"E9E9EAEAEAEBEBECECEDEDEEEEEFEFF0F0F1F1F1F2F2F3F3F4F4F5F5F6F6F7F7";
constant INIT_H_TH0_75 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH0_75 : bit_vector(255 downto 0) := X"DADADBDBDCDCDDDDDEDEDEDFDFE0E0E1E1E2E2E3E3E4E4E4E5E5E6E6E7E7E8E8";
constant INIT_H_TH0_76 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH0_76 : bit_vector(255 downto 0) := X"CBCCCCCDCDCECECECFCFD0D0D1D1D2D2D3D3D3D4D4D5D5D6D6D7D7D8D8D9D9D9";
constant INIT_H_TH0_77 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH0_77 : bit_vector(255 downto 0) := X"BDBDBEBEBFBFC0C0C0C1C1C2C2C3C3C4C4C4C5C5C6C6C7C7C8C8C9C9C9CACACB";
constant INIT_H_TH0_78 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH0_78 : bit_vector(255 downto 0) := X"AEAFAFB0B0B1B1B2B2B3B3B3B4B4B5B5B6B6B7B7B7B8B8B9B9BABABBBBBBBCBC";
constant INIT_H_TH0_79 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH0_79 : bit_vector(255 downto 0) := X"A0A1A1A2A2A2A3A3A4A4A5A5A6A6A6A7A7A8A8A9A9AAAAAAABABACACADADAEAE";
constant INIT_H_TH0_7A : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH0_7A : bit_vector(255 downto 0) := X"92939394949495959696979797989899999A9A9B9B9B9C9C9D9D9E9E9F9F9FA0";
constant INIT_H_TH0_7B : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH0_7B : bit_vector(255 downto 0) := X"848585868686878788888989898A8A8B8B8C8C8D8D8D8E8E8F8F909090919192";
constant INIT_H_TH0_7C : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH0_7C : bit_vector(255 downto 0) := X"76777778787979797A7A7B7B7C7C7C7D7D7E7E7F7F8080808181828283838384";
constant INIT_H_TH0_7D : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH0_7D : bit_vector(255 downto 0) := X"69696A6A6A6B6B6C6C6D6D6D6E6E6F6F70707071717272737373747475757676";
constant INIT_H_TH0_7E : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH0_7E : bit_vector(255 downto 0) := X"5B5C5C5C5D5D5E5E5F5F5F606061616262626363646465656566666767676868";
constant INIT_H_TH0_7F : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH0_7F : bit_vector(255 downto 0) := X"4E4E4F4F4F5050515152525253535454545555565657575758585959595A5A5B";
constant INIT_H_TH1_00 : bit_vector(255 downto 0) := X"2626262626262626262626262626262626262626262626262626262626262626";
constant INIT_L_TH1_00 : bit_vector(255 downto 0) := X"016FE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1";
constant INIT_H_TH1_01 : bit_vector(255 downto 0) := X"1D1D1D1D1E1E1E1E1E1F1F1F1F20202020212121212222222323232424242525";
constant INIT_L_TH1_01 : bit_vector(255 downto 0) := X"4070A1D306396EA4DB134C87C3003F7FC1044A90D92471C01165BB1470D03298";
constant INIT_H_TH1_02 : bit_vector(255 downto 0) := X"1818181819191919191919191A1A1A1A1A1A1A1B1B1B1B1B1B1C1C1C1C1C1C1D";
constant INIT_L_TH1_02 : bit_vector(255 downto 0) := X"98B6D4F21131507091B2D3F5183B5E82A6CBF1173D648CB5DE07325D89B5E311";
constant INIT_H_TH1_03 : bit_vector(255 downto 0) := X"1515151515151516161616161616161616161717171717171717171818181818";
constant INIT_L_TH1_03 : bit_vector(255 downto 0) := X"788DA3B8CEE4FB11283F566E859DB5CEE7FF19324C66809BB5D1EC0824405D7A";
constant INIT_H_TH1_04 : bit_vector(255 downto 0) := X"1313131313131313131313131314141414141414141414141414141515151515";
constant INIT_L_TH1_04 : bit_vector(255 downto 0) := X"2334445566778899ABBCCEDFF10316283A4D60738699ACC0D4E8FC1024394E63";
constant INIT_H_TH1_05 : bit_vector(255 downto 0) := X"1111111111111111111111111111121212121212121212121212121212121313";
constant INIT_L_TH1_05 : bit_vector(255 downto 0) := X"4B586673818E9CAAB8C6D4E2F1FF0D1C2B39485766758594A4B3C3D3E3F30313";
constant INIT_H_TH1_06 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F1010101010101010101010101010101010101010101111111111";
constant INIT_L_TH1_06 : bit_vector(255 downto 0) := X"C5D0DCE7F2FE0915202C38434F5B67737F8C98A4B0BDC9D6E3EFFC091623303E";
constant INIT_H_TH1_07 : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_TH1_07 : bit_vector(255 downto 0) := X"7B848E98A1ABB5BFC9D3DDE7F1FB050F1A242E39434E58636E78838E99A4AFBA";
constant INIT_H_TH1_08 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_TH1_08 : bit_vector(255 downto 0) := X"5C656D767E878F98A0A9B2BAC3CCD5DEE7F0F9020B141D262F39424B555E6871";
constant INIT_H_TH1_09 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_TH1_09 : bit_vector(255 downto 0) := X"60686F777E868D959DA4ACB4BBC3CBD3DBE2EAF2FA020A121A232B333B434C54";
constant INIT_H_TH1_0A : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_TH1_0A : bit_vector(255 downto 0) := X"80868D949AA1A8AFB6BCC3CAD1D8DFE6EDF4FB020910171F262D343C434A5259";
constant INIT_H_TH1_0B : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_TH1_0B : bit_vector(255 downto 0) := X"B5BBC1C7CDD3DAE0E6ECF2F8FF050B11181E242B31383E454B52585F656C7279";
constant INIT_H_TH1_0C : bit_vector(255 downto 0) := X"090A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_TH1_0C : bit_vector(255 downto 0) := X"FD02080D13191E24292F353A40464B51575D62686E747A7F858B91979DA3A9AF";
constant INIT_H_TH1_0D : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_TH1_0D : bit_vector(255 downto 0) := X"54595E63686E73787D82878C92979CA1A7ACB1B7BCC1C7CCD1D7DCE1E7ECF2F7";
constant INIT_H_TH1_0E : bit_vector(255 downto 0) := X"0808080808080808080808080808080909090909090909090909090909090909";
constant INIT_L_TH1_0E : bit_vector(255 downto 0) := X"B9BDC2C7CBD0D5DADEE3E8EDF1F6FB00050A0F13181D22272C31363B40454A4F";
constant INIT_H_TH1_0F : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_TH1_0F : bit_vector(255 downto 0) := X"282D31353A3E43474B5054595D62666B6F74787D81868A8F93989DA1A6ABAFB4";
constant INIT_H_TH1_10 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707080808080808080808";
constant INIT_L_TH1_10 : bit_vector(255 downto 0) := X"A2A6AAAEB2B6BBBFC3C7CBCFD3D7DCE0E4E8ECF1F5F9FD02060A0E13171B2024";
constant INIT_H_TH1_11 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_TH1_11 : bit_vector(255 downto 0) := X"24282C3034383B3F43474B4F53565A5E62666A6E72767A7E82868A8E92969A9E";
constant INIT_H_TH1_12 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606070707070707070707";
constant INIT_L_TH1_12 : bit_vector(255 downto 0) := X"AEB2B6B9BDC0C4C8CBCFD3D6DADEE1E5E9ECF0F4F7FBFF03060A0E1215191D21";
constant INIT_H_TH1_13 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_TH1_13 : bit_vector(255 downto 0) := X"3F43464A4D5054575B5E6165686C6F73767A7D8184888B8F9296999DA0A4A7AB";
constant INIT_H_TH1_14 : bit_vector(255 downto 0) := X"0505050505050505050505050506060606060606060606060606060606060606";
constant INIT_L_TH1_14 : bit_vector(255 downto 0) := X"D6DADDE0E3E6EAEDF0F3F7FAFD0004070A0D1114171B1E2125282B2F3235393C";
constant INIT_H_TH1_15 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_TH1_15 : bit_vector(255 downto 0) := X"7376797C7F8285888B8E9195989B9EA1A4A7AAADB0B4B7BABDC0C3C6CACDD0D3";
constant INIT_H_TH1_16 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_TH1_16 : bit_vector(255 downto 0) := X"14171A1D202326292C2F3134373A3D404346494C4F5255585B5E6164676A6D70";
constant INIT_H_TH1_17 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040405050505050505";
constant INIT_L_TH1_17 : bit_vector(255 downto 0) := X"BBBDC0C3C6C8CBCED1D3D6D9DCDFE1E4E7EAEDEFF2F5F8FBFE000306090C0F12";
constant INIT_H_TH1_18 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_TH1_18 : bit_vector(255 downto 0) := X"65676A6D6F7275777A7C7F8284878A8C8F9295979A9D9FA2A5A7AAADB0B2B5B8";
constant INIT_H_TH1_19 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_TH1_19 : bit_vector(255 downto 0) := X"1315181A1D1F222427292C2F313436393B3E404346484B4D505255585A5D5F62";
constant INIT_H_TH1_1A : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030304040404040404";
constant INIT_L_TH1_1A : bit_vector(255 downto 0) := X"C4C7C9CBCED0D3D5D8DADCDFE1E4E6E9EBEEF0F2F5F7FAFCFF010406090B0E10";
constant INIT_H_TH1_1B : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_TH1_1B : bit_vector(255 downto 0) := X"797B7E80828587898B8E909295979A9C9EA1A3A5A8AAACAFB1B3B6B8BBBDBFC2";
constant INIT_H_TH1_1C : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_TH1_1C : bit_vector(255 downto 0) := X"313335373A3C3E40424547494B4E50525457595B5D60626467696B6D70727477";
constant INIT_H_TH1_1D : bit_vector(255 downto 0) := X"0202020202020202020203030303030303030303030303030303030303030303";
constant INIT_L_TH1_1D : bit_vector(255 downto 0) := X"EBEDEFF2F4F6F8FAFCFE01030507090B0E10121416181B1D1F212326282A2C2E";
constant INIT_H_TH1_1E : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_TH1_1E : bit_vector(255 downto 0) := X"A8AAACAEB0B2B4B7B9BBBDBFC1C3C5C7C9CBCDD0D2D4D6D8DADCDEE0E3E5E7E9";
constant INIT_H_TH1_1F : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_TH1_1F : bit_vector(255 downto 0) := X"686A6C6D6F71737577797B7D7F818486888A8C8E90929496989A9C9EA0A2A4A6";
constant INIT_H_TH1_20 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_TH1_20 : bit_vector(255 downto 0) := X"292B2D2F31333537393B3C3E40424446484A4C4E50525456585A5C5E60626466";
constant INIT_H_TH1_21 : bit_vector(255 downto 0) := X"0101010101010101010102020202020202020202020202020202020202020202";
constant INIT_L_TH1_21 : bit_vector(255 downto 0) := X"EDEFF1F3F4F6F8FAFCFE0001030507090B0D0F10121416181A1C1E2022232527";
constant INIT_H_TH1_22 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_TH1_22 : bit_vector(255 downto 0) := X"B3B4B6B8BABCBDBFC1C3C5C6C8CACCCED0D1D3D5D7D9DBDCDEE0E2E4E6E7E9EB";
constant INIT_H_TH1_23 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_TH1_23 : bit_vector(255 downto 0) := X"7A7C7E7F81838586888A8C8D8F91939496989A9C9D9FA1A3A4A6A8AAACADAFB1";
constant INIT_H_TH1_24 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_TH1_24 : bit_vector(255 downto 0) := X"444547494A4C4E4F51535456585A5B5D5F6062646667696B6C6E707273757778";
constant INIT_H_TH1_25 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_TH1_25 : bit_vector(255 downto 0) := X"0E1012131517181A1C1D1F2122242527292A2C2E2F3133343638393B3D3E4042";
constant INIT_H_TH1_26 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000010101010101010101";
constant INIT_L_TH1_26 : bit_vector(255 downto 0) := X"DBDDDEE0E1E3E5E6E8E9EBEDEEF0F1F3F5F6F8F9FBFDFE0001030506080A0B0D";
constant INIT_H_TH1_27 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_TH1_27 : bit_vector(255 downto 0) := X"A9AAACAEAFB1B2B4B5B7B8BABCBDBFC0C2C3C5C6C8CACBCDCED0D1D3D5D6D8D9";
constant INIT_H_TH1_28 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_TH1_28 : bit_vector(255 downto 0) := X"787A7B7D7E808183848687898A8C8D8F9092939597989A9B9D9EA0A1A3A4A6A7";
constant INIT_H_TH1_29 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_TH1_29 : bit_vector(255 downto 0) := X"494A4C4D4F505253555658595B5C5E5F606263656668696B6C6E6F7172747577";
constant INIT_H_TH1_2A : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_TH1_2A : bit_vector(255 downto 0) := X"1B1C1E1F212223252628292B2C2D2F303233353638393A3C3D3F404243454648";
constant INIT_H_TH1_2B : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000";
constant INIT_L_TH1_2B : bit_vector(255 downto 0) := X"EEEFF1F2F4F5F6F8F9FBFCFDFF000103040607090A0B0D0E1011121415171819";
constant INIT_H_TH1_2C : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_TH1_2C : bit_vector(255 downto 0) := X"C2C4C5C6C8C9CACCCDCED0D1D3D4D5D7D8D9DBDCDDDFE0E2E3E4E6E7E8EAEBED";
constant INIT_H_TH1_2D : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_TH1_2D : bit_vector(255 downto 0) := X"98999A9C9D9E9FA1A2A3A5A6A7A9AAABADAEAFB1B2B3B5B6B7B9BABCBDBEC0C1";
constant INIT_H_TH1_2E : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_TH1_2E : bit_vector(255 downto 0) := X"6E6F707273747677787A7B7C7D7F80818384858788898A8C8D8E909192949596";
constant INIT_H_TH1_2F : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_TH1_2F : bit_vector(255 downto 0) := X"454748494A4C4D4E4F51525354565758595B5C5D5F60616264656668696A6B6D";
constant INIT_H_TH1_30 : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_TH1_30 : bit_vector(255 downto 0) := X"1E1F20212224252627292A2B2C2E2F30313334353638393A3B3C3E3F40424344";
constant INIT_H_TH1_31 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_TH1_31 : bit_vector(255 downto 0) := X"F7F8F9FAFCFDFEFF00020304050608090A0B0C0E0F10111314151617191A1B1C";
constant INIT_H_TH1_32 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH1_32 : bit_vector(255 downto 0) := X"D1D2D3D4D5D7D8D9DADBDDDEDFE0E1E2E4E5E6E7E8EAEBECEDEEF0F1F2F3F4F6";
constant INIT_H_TH1_33 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH1_33 : bit_vector(255 downto 0) := X"ACADAEAFB0B1B3B4B5B6B7B8B9BBBCBDBEBFC0C2C3C4C5C6C7C9CACBCCCDCED0";
constant INIT_H_TH1_34 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH1_34 : bit_vector(255 downto 0) := X"87888A8B8C8D8E8F9091939495969798999B9C9D9E9FA0A1A2A4A5A6A7A8A9AB";
constant INIT_H_TH1_35 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH1_35 : bit_vector(255 downto 0) := X"6465666768696A6B6D6E6F7071727374757778797A7B7C7D7E7F818283848586";
constant INIT_H_TH1_36 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH1_36 : bit_vector(255 downto 0) := X"41424344454647484A4B4C4D4E4F5051525354565758595A5B5C5D5E5F606263";
constant INIT_H_TH1_37 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH1_37 : bit_vector(255 downto 0) := X"1F202122232425262728292A2B2D2E2F303132333435363738393A3C3D3E3F40";
constant INIT_H_TH1_38 : bit_vector(255 downto 0) := X"FDFDFDFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_TH1_38 : bit_vector(255 downto 0) := X"FDFEFF0001030405060708090A0B0C0D0E0F1011121314151617181A1B1C1D1E";
constant INIT_H_TH1_39 : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH1_39 : bit_vector(255 downto 0) := X"DDDEDFE0E1E2E3E4E5E6E7E8E9EAEBECEDEEEFF0F1F2F3F4F5F6F7F8F9FAFBFC";
constant INIT_H_TH1_3A : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH1_3A : bit_vector(255 downto 0) := X"BCBDBEBFC0C1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADB";
constant INIT_H_TH1_3B : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH1_3B : bit_vector(255 downto 0) := X"9D9E9FA0A1A2A3A4A5A6A7A8A9AAABABACADAEAFB0B1B2B3B4B5B6B7B8B9BABB";
constant INIT_H_TH1_3C : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH1_3C : bit_vector(255 downto 0) := X"7E7F80818283848585868788898A8B8C8D8E8F909192939495969798999A9B9C";
constant INIT_H_TH1_3D : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH1_3D : bit_vector(255 downto 0) := X"5F606162636465666768696A6B6C6D6E6F6F707172737475767778797A7B7C7D";
constant INIT_H_TH1_3E : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH1_3E : bit_vector(255 downto 0) := X"4142434445464748494A4B4C4D4E4E4F505152535455565758595A5B5C5D5D5E";
constant INIT_H_TH1_3F : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH1_3F : bit_vector(255 downto 0) := X"2425262728292A2B2B2C2D2E2F30313233343536363738393A3B3C3D3E3F4041";
constant INIT_H_TH1_40 : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_TH1_40 : bit_vector(255 downto 0) := X"0708090A0B0C0D0E0E0F10111213141516171718191A1B1C1D1E1F2021212223";
constant INIT_H_TH1_41 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFDFDFDFDFDFDFDFD";
constant INIT_L_TH1_41 : bit_vector(255 downto 0) := X"EBECEDEEEEEFF0F1F2F3F4F5F6F6F7F8F9FAFBFCFDFEFEFF0001020304050606";
constant INIT_H_TH1_42 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH1_42 : bit_vector(255 downto 0) := X"CFD0D1D2D3D3D4D5D6D7D8D9D9DADBDCDDDEDFE0E0E1E2E3E4E5E6E7E7E8E9EA";
constant INIT_H_TH1_43 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH1_43 : bit_vector(255 downto 0) := X"B4B5B5B6B7B8B9BABBBBBCBDBEBFC0C0C1C2C3C4C5C6C6C7C8C9CACBCCCDCDCE";
constant INIT_H_TH1_44 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH1_44 : bit_vector(255 downto 0) := X"999A9A9B9C9D9E9F9FA0A1A2A3A4A4A5A6A7A8A9AAAAABACADAEAFAFB0B1B2B3";
constant INIT_H_TH1_45 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH1_45 : bit_vector(255 downto 0) := X"7E7F8081828283848586868788898A8B8B8C8D8E8F9090919293949595969798";
constant INIT_H_TH1_46 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH1_46 : bit_vector(255 downto 0) := X"646566676768696A6B6B6C6D6E6F6F7071727374747576777878797A7B7C7D7D";
constant INIT_H_TH1_47 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH1_47 : bit_vector(255 downto 0) := X"4A4B4C4D4E4E4F5051525253545556565758595A5A5B5C5D5E5E5F6061626363";
constant INIT_H_TH1_48 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH1_48 : bit_vector(255 downto 0) := X"31323333343536373738393A3B3B3C3D3E3F3F4041424243444546464748494A";
constant INIT_H_TH1_49 : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH1_49 : bit_vector(255 downto 0) := X"18191A1B1B1C1D1E1E1F202122222324252526272829292A2B2C2C2D2E2F3030";
constant INIT_H_TH1_4A : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_TH1_4A : bit_vector(255 downto 0) := X"000001020303040506070708090A0A0B0C0D0D0E0F1011111213141415161717";
constant INIT_H_TH1_4B : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH1_4B : bit_vector(255 downto 0) := X"E8E8E9EAEBEBECEDEEEEEFF0F1F1F2F3F4F4F5F6F7F7F8F9FAFAFBFCFDFDFEFF";
constant INIT_H_TH1_4C : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH1_4C : bit_vector(255 downto 0) := X"D0D0D1D2D3D3D4D5D6D6D7D8D9D9DADBDCDCDDDEDFDFE0E1E2E2E3E4E5E5E6E7";
constant INIT_H_TH1_4D : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH1_4D : bit_vector(255 downto 0) := X"B8B9BABABBBCBDBDBEBFC0C0C1C2C2C3C4C5C5C6C7C8C8C9CACBCBCCCDCDCECF";
constant INIT_H_TH1_4E : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH1_4E : bit_vector(255 downto 0) := X"A1A2A3A3A4A5A5A6A7A8A8A9AAAAABACADADAEAFB0B0B1B2B2B3B4B5B5B6B7B7";
constant INIT_H_TH1_4F : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH1_4F : bit_vector(255 downto 0) := X"8A8B8C8C8D8E8F8F90919192939494959696979898999A9B9B9C9D9E9E9FA0A0";
constant INIT_H_TH1_50 : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH1_50 : bit_vector(255 downto 0) := X"7474757677777879797A7B7B7C7D7E7E7F80808182838384858586878788898A";
constant INIT_H_TH1_51 : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH1_51 : bit_vector(255 downto 0) := X"5E5E5F6060616262636464656667676869696A6B6B6C6D6E6E6F707071727273";
constant INIT_H_TH1_52 : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH1_52 : bit_vector(255 downto 0) := X"4848494A4A4B4C4C4D4E4F4F5051515253535455555657575859595A5B5C5C5D";
constant INIT_H_TH1_53 : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH1_53 : bit_vector(255 downto 0) := X"32333334353536373738393A3A3B3C3C3D3E3E3F404041424243444445464647";
constant INIT_H_TH1_54 : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH1_54 : bit_vector(255 downto 0) := X"1D1D1E1F1F2021212223232425252627272829292A2B2B2C2D2D2E2F2F303131";
constant INIT_H_TH1_55 : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH1_55 : bit_vector(255 downto 0) := X"0808090A0A0B0C0C0D0E0E0F1010111212131414151616171818191A1A1B1B1C";
constant INIT_H_TH1_56 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_TH1_56 : bit_vector(255 downto 0) := X"F3F4F4F5F6F6F7F8F8F9F9FAFBFBFCFDFDFEFFFF000101020303040505060607";
constant INIT_H_TH1_57 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_57 : bit_vector(255 downto 0) := X"DFDFE0E0E1E2E2E3E4E4E5E6E6E7E7E8E9E9EAEBEBECEDEDEEEFEFF0F0F1F2F2";
constant INIT_H_TH1_58 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_58 : bit_vector(255 downto 0) := X"CACBCCCCCDCDCECFCFD0D1D1D2D2D3D4D4D5D6D6D7D8D8D9D9DADBDBDCDDDDDE";
constant INIT_H_TH1_59 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_59 : bit_vector(255 downto 0) := X"B6B7B8B8B9B9BABBBBBCBDBDBEBEBFC0C0C1C2C2C3C3C4C5C5C6C7C7C8C8C9CA";
constant INIT_H_TH1_5A : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_5A : bit_vector(255 downto 0) := X"A3A3A4A4A5A6A6A7A7A8A9A9AAABABACACADAEAEAFB0B0B1B1B2B3B3B4B4B5B6";
constant INIT_H_TH1_5B : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_5B : bit_vector(255 downto 0) := X"8F90909192929393949595969697989899999A9B9B9C9C9D9E9E9FA0A0A1A1A2";
constant INIT_H_TH1_5C : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_5C : bit_vector(255 downto 0) := X"7C7C7D7E7E7F7F808181828283848485858687878888898A8A8B8B8C8D8D8E8E";
constant INIT_H_TH1_5D : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_5D : bit_vector(255 downto 0) := X"69696A6B6B6C6C6D6E6E6F6F70717172727373747575767677787879797A7B7B";
constant INIT_H_TH1_5E : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_5E : bit_vector(255 downto 0) := X"5657575858595A5A5B5B5C5C5D5E5E5F5F606161626263636465656666676868";
constant INIT_H_TH1_5F : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_5F : bit_vector(255 downto 0) := X"43444545464647474849494A4A4B4C4C4D4D4E4E4F5050515152535354545555";
constant INIT_H_TH1_60 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_60 : bit_vector(255 downto 0) := X"3132323333343435363637373838393A3A3B3B3C3D3D3E3E3F3F404141424243";
constant INIT_H_TH1_61 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_61 : bit_vector(255 downto 0) := X"1F1F20212122222323242525262627272829292A2A2B2B2C2C2D2E2E2F2F3030";
constant INIT_H_TH1_62 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_62 : bit_vector(255 downto 0) := X"0D0E0E0F0F1010111112131314141515161617181819191A1A1B1C1C1D1D1E1E";
constant INIT_H_TH1_63 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_TH1_63 : bit_vector(255 downto 0) := X"FBFCFCFDFDFEFFFF0000010102020303040505060607070808090A0A0B0B0C0C";
constant INIT_H_TH1_64 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_64 : bit_vector(255 downto 0) := X"EAEAEBEBECECEDEDEEEFEFF0F0F1F1F2F2F3F3F4F5F5F6F6F7F7F8F8F9FAFAFB";
constant INIT_H_TH1_65 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_65 : bit_vector(255 downto 0) := X"D8D9D9DADADBDCDCDDDDDEDEDFDFE0E0E1E1E2E3E3E4E4E5E5E6E6E7E7E8E9E9";
constant INIT_H_TH1_66 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_66 : bit_vector(255 downto 0) := X"C7C8C8C9C9CACACBCBCCCCCDCECECFCFD0D0D1D1D2D2D3D3D4D5D5D6D6D7D7D8";
constant INIT_H_TH1_67 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_67 : bit_vector(255 downto 0) := X"B6B7B7B8B8B9B9BABABBBBBCBCBDBEBEBFBFC0C0C1C1C2C2C3C3C4C4C5C6C6C7";
constant INIT_H_TH1_68 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_68 : bit_vector(255 downto 0) := X"A5A6A6A7A7A8A8A9AAAAABABACACADADAEAEAFAFB0B0B1B1B2B2B3B3B4B5B5B6";
constant INIT_H_TH1_69 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_69 : bit_vector(255 downto 0) := X"959596969797989899999A9A9B9B9C9C9D9E9E9F9FA0A0A1A1A2A2A3A3A4A4A5";
constant INIT_H_TH1_6A : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_6A : bit_vector(255 downto 0) := X"84858586868787888889898A8A8B8B8C8C8D8D8E8F8F90909191929293939494";
constant INIT_H_TH1_6B : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_6B : bit_vector(255 downto 0) := X"74747575767777787879797A7A7B7B7C7C7D7D7E7E7F7F808081818282838384";
constant INIT_H_TH1_6C : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_6C : bit_vector(255 downto 0) := X"6464656566666767686869696A6A6B6B6C6C6D6D6E6E6F6F7070717172727373";
constant INIT_H_TH1_6D : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_6D : bit_vector(255 downto 0) := X"5454555556565757585859595A5A5B5B5C5C5D5D5E5E5F5F6060616162626363";
constant INIT_H_TH1_6E : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_6E : bit_vector(255 downto 0) := X"44454546464747484849494A4A4B4B4C4C4C4D4D4E4E4F4F5050515152525353";
constant INIT_H_TH1_6F : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_6F : bit_vector(255 downto 0) := X"35353536363737383839393A3A3B3B3C3C3D3D3E3E3F3F404041414242434344";
constant INIT_H_TH1_70 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_70 : bit_vector(255 downto 0) := X"252626262727282829292A2A2B2B2C2C2D2D2E2E2F2F30303131323233333434";
constant INIT_H_TH1_71 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_71 : bit_vector(255 downto 0) := X"16161717181819191A1A1A1B1B1C1C1D1D1E1E1F1F2020212122222323242425";
constant INIT_H_TH1_72 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_72 : bit_vector(255 downto 0) := X"070707080809090A0A0B0B0C0C0D0D0E0E0F0F10101011111212131314141515";
constant INIT_H_TH1_73 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_TH1_73 : bit_vector(255 downto 0) := X"F8F8F8F9F9FAFAFBFBFCFCFDFDFEFEFFFFFF0000010102020303040405050606";
constant INIT_H_TH1_74 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH1_74 : bit_vector(255 downto 0) := X"E9E9EAEAEAEBEBECECEDEDEEEEEFEFF0F0F1F1F1F2F2F3F3F4F4F5F5F6F6F7F7";
constant INIT_H_TH1_75 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH1_75 : bit_vector(255 downto 0) := X"DADADBDBDCDCDDDDDEDEDEDFDFE0E0E1E1E2E2E3E3E4E4E4E5E5E6E6E7E7E8E8";
constant INIT_H_TH1_76 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH1_76 : bit_vector(255 downto 0) := X"CBCCCCCDCDCECECECFCFD0D0D1D1D2D2D3D3D3D4D4D5D5D6D6D7D7D8D8D9D9D9";
constant INIT_H_TH1_77 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH1_77 : bit_vector(255 downto 0) := X"BDBDBEBEBFBFC0C0C0C1C1C2C2C3C3C4C4C4C5C5C6C6C7C7C8C8C9C9C9CACACB";
constant INIT_H_TH1_78 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH1_78 : bit_vector(255 downto 0) := X"AEAFAFB0B0B1B1B2B2B3B3B3B4B4B5B5B6B6B7B7B7B8B8B9B9BABABBBBBBBCBC";
constant INIT_H_TH1_79 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH1_79 : bit_vector(255 downto 0) := X"A0A1A1A2A2A2A3A3A4A4A5A5A6A6A6A7A7A8A8A9A9AAAAAAABABACACADADAEAE";
constant INIT_H_TH1_7A : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH1_7A : bit_vector(255 downto 0) := X"92939394949495959696979797989899999A9A9B9B9B9C9C9D9D9E9E9F9F9FA0";
constant INIT_H_TH1_7B : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH1_7B : bit_vector(255 downto 0) := X"848585868686878788888989898A8A8B8B8C8C8D8D8D8E8E8F8F909090919192";
constant INIT_H_TH1_7C : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH1_7C : bit_vector(255 downto 0) := X"76777778787979797A7A7B7B7C7C7C7D7D7E7E7F7F8080808181828283838384";
constant INIT_H_TH1_7D : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH1_7D : bit_vector(255 downto 0) := X"69696A6A6A6B6B6C6C6D6D6D6E6E6F6F70707071717272737373747475757676";
constant INIT_H_TH1_7E : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH1_7E : bit_vector(255 downto 0) := X"5B5C5C5C5D5D5E5E5F5F5F606061616262626363646465656566666767676868";
constant INIT_H_TH1_7F : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_TH1_7F : bit_vector(255 downto 0) := X"4E4E4F4F4F5050515152525253535454545555565657575758585959595A5A5B";
constant INIT_H_HUM_00 : bit_vector(255 downto 0) := X"F7F7F7F7F7F7F7F7F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6";
constant INIT_L_HUM_00 : bit_vector(255 downto 0) := X"1814110E0B080401FEFBF8F4F1EEEBE8E4E1DEDBD8D4D1CECBC8C4C1BEBBB8B4";
constant INIT_H_HUM_01 : bit_vector(255 downto 0) := X"F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7";
constant INIT_L_HUM_01 : bit_vector(255 downto 0) := X"7E7B7874716E6B6864615E5B5854514E4B4844413E3B3834312E2B2824211E1B";
constant INIT_H_HUM_02 : bit_vector(255 downto 0) := X"F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7";
constant INIT_L_HUM_02 : bit_vector(255 downto 0) := X"E4E1DEDBD8D4D1CECBC8C4C1BEBBB8B4B1AEABA8A4A19E9B9894918E8B888481";
constant INIT_H_HUM_03 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F7F7F7F7F7F7F7F7";
constant INIT_L_HUM_03 : bit_vector(255 downto 0) := X"4B4844413E3B3834312E2B2824211E1B1814110E0B080401FEFBF8F4F1EEEBE8";
constant INIT_H_HUM_04 : bit_vector(255 downto 0) := X"F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_HUM_04 : bit_vector(255 downto 0) := X"B1AEABA8A4A19E9B9894918E8B8884817E7B7874716E6B6864615E5B5854514E";
constant INIT_H_HUM_05 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8";
constant INIT_L_HUM_05 : bit_vector(255 downto 0) := X"1814110E0B080401FEFBF8F4F1EEEBE8E4E1DEDBD8D4D1CECBC8C4C1BEBBB8B4";
constant INIT_H_HUM_06 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_HUM_06 : bit_vector(255 downto 0) := X"7E7B7874716E6B6864615E5B5854514E4B4844413E3B3834312E2B2824211E1B";
constant INIT_H_HUM_07 : bit_vector(255 downto 0) := X"F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9";
constant INIT_L_HUM_07 : bit_vector(255 downto 0) := X"E4E1DEDBD8D4D1CECBC8C4C1BEBBB8B4B1AEABA8A4A19E9B9894918E8B888481";
constant INIT_H_HUM_08 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAF9F9F9F9F9F9F9F9";
constant INIT_L_HUM_08 : bit_vector(255 downto 0) := X"4B4844413E3B3834312E2B2824211E1B1814110E0B080401FEFBF8F4F1EEEBE8";
constant INIT_H_HUM_09 : bit_vector(255 downto 0) := X"FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_HUM_09 : bit_vector(255 downto 0) := X"B1AEABA8A4A19E9B9894918E8B8884817E7B7874716E6B6864615E5B5854514E";
constant INIT_H_HUM_0A : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA";
constant INIT_L_HUM_0A : bit_vector(255 downto 0) := X"1814110E0B080401FEFBF8F4F1EEEBE8E4E1DEDBD8D4D1CECBC8C4C1BEBBB8B4";
constant INIT_H_HUM_0B : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_HUM_0B : bit_vector(255 downto 0) := X"7E7B7874716E6B6864615E5B5854514E4B4844413E3B3834312E2B2824211E1B";
constant INIT_H_HUM_0C : bit_vector(255 downto 0) := X"FBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB";
constant INIT_L_HUM_0C : bit_vector(255 downto 0) := X"E4E1DEDBD8D4D1CECBC8C4C1BEBBB8B4B1AEABA8A4A19E9B9894918E8B888481";
constant INIT_H_HUM_0D : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFBFBFBFBFBFBFBFB";
constant INIT_L_HUM_0D : bit_vector(255 downto 0) := X"4B4844413E3B3834312E2B2824211E1B1814110E0B080401FEFBF8F4F1EEEBE8";
constant INIT_H_HUM_0E : bit_vector(255 downto 0) := X"FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_HUM_0E : bit_vector(255 downto 0) := X"B1AEABA8A4A19E9B9894918E8B8884817E7B7874716E6B6864615E5B5854514E";
constant INIT_H_HUM_0F : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC";
constant INIT_L_HUM_0F : bit_vector(255 downto 0) := X"1814110E0B080401FEFBF8F4F1EEEBE8E4E1DEDBD8D4D1CECBC8C4C1BEBBB8B4";
constant INIT_H_HUM_10 : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_HUM_10 : bit_vector(255 downto 0) := X"7E7B7874716E6B6864615E5B5854514E4B4844413E3B3834312E2B2824211E1B";
constant INIT_H_HUM_11 : bit_vector(255 downto 0) := X"FDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD";
constant INIT_L_HUM_11 : bit_vector(255 downto 0) := X"E4E1DEDBD8D4D1CECBC8C4C1BEBBB8B4B1AEABA8A4A19E9B9894918E8B888481";
constant INIT_H_HUM_12 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFDFDFDFDFDFDFDFD";
constant INIT_L_HUM_12 : bit_vector(255 downto 0) := X"4B4844413E3B3834312E2B2824211E1B1814110E0B080401FEFBF8F4F1EEEBE8";
constant INIT_H_HUM_13 : bit_vector(255 downto 0) := X"FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_HUM_13 : bit_vector(255 downto 0) := X"B1AEABA8A4A19E9B9894918E8B8884817E7B7874716E6B6864615E5B5854514E";
constant INIT_H_HUM_14 : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE";
constant INIT_L_HUM_14 : bit_vector(255 downto 0) := X"1714110E0B070401FEFBF7F4F1EEEBE7E4E1DEDBD7D4D1CECBC7C4C1BEBBB8B4";
constant INIT_H_HUM_15 : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_HUM_15 : bit_vector(255 downto 0) := X"7E7B7774716E6B6764615E5B5754514E4B4744413E3B3734312E2B2724211E1B";
constant INIT_H_HUM_16 : bit_vector(255 downto 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant INIT_L_HUM_16 : bit_vector(255 downto 0) := X"E4E1DEDBD7D4D1CECBC7C4C1BEBBB7B4B1AEABA7A4A19E9B9794918E8B878481";
constant INIT_H_HUM_17 : bit_vector(255 downto 0) := X"000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFF";
constant INIT_L_HUM_17 : bit_vector(255 downto 0) := X"4A4643403D3A3633302D2A2623201D1A1613100D0A060300FEFBF7F4F1EEEBE7";
constant INIT_H_HUM_18 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_HUM_18 : bit_vector(255 downto 0) := X"B0ADAAA6A3A09D9A9693908D8A8683807D7A7673706D6A6663605D5A5653504D";
constant INIT_H_HUM_19 : bit_vector(255 downto 0) := X"0101010101010101000000000000000000000000000000000000000000000000";
constant INIT_L_HUM_19 : bit_vector(255 downto 0) := X"1613100D0A060300FDFAF6F3F0EDEAE6E3E0DDDAD6D3D0CDCAC6C3C0BDBAB6B3";
constant INIT_H_HUM_1A : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_HUM_1A : bit_vector(255 downto 0) := X"7D7A7673706D6A6663605D5A5653504D4A4643403D3A3633302D2A2623201D1A";
constant INIT_H_HUM_1B : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_HUM_1B : bit_vector(255 downto 0) := X"E3E0DDDAD6D3D0CDCAC6C3C0BDBAB6B3B0ADAAA6A3A09D9A9693908D8A868380";
constant INIT_H_HUM_1C : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020101010101010101";
constant INIT_L_HUM_1C : bit_vector(255 downto 0) := X"4A4643403D3A3633302D2A2623201D1A1613100D0A060300FDFAF6F3F0EDEAE6";
constant INIT_H_HUM_1D : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_HUM_1D : bit_vector(255 downto 0) := X"B0ADAAA6A3A09D9A9693908D8A8683807D7A7673706D6A6663605D5A5653504D";
constant INIT_H_HUM_1E : bit_vector(255 downto 0) := X"0303030303030303020202020202020202020202020202020202020202020202";
constant INIT_L_HUM_1E : bit_vector(255 downto 0) := X"1613100D0A060300FDFAF6F3F0EDEAE6E3E0DDDAD6D3D0CDCAC6C3C0BDBAB6B3";
constant INIT_H_HUM_1F : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_HUM_1F : bit_vector(255 downto 0) := X"7D7A7673706D6A6663605D5A5653504D4A4643403D3A3633302D2A2623201D1A";
constant INIT_H_HUM_20 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_HUM_20 : bit_vector(255 downto 0) := X"E3E0DDDAD6D3D0CDCAC6C3C0BDBAB6B3B0ADAAA6A3A09D9A9693908D8A868380";
constant INIT_H_HUM_21 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040303030303030303";
constant INIT_L_HUM_21 : bit_vector(255 downto 0) := X"4A4643403D3A3633302D2A2623201D1A1613100D0A060300FDFAF6F3F0EDEAE6";
constant INIT_H_HUM_22 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_HUM_22 : bit_vector(255 downto 0) := X"B0ADAAA6A3A09D9A9693908D8A8683807D7A7673706D6A6663605D5A5653504D";
constant INIT_H_HUM_23 : bit_vector(255 downto 0) := X"0505050505050505040404040404040404040404040404040404040404040404";
constant INIT_L_HUM_23 : bit_vector(255 downto 0) := X"1613100D0A060300FDFAF6F3F0EDEAE6E3E0DDDAD6D3D0CDCAC6C3C0BDBAB6B3";
constant INIT_H_HUM_24 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_HUM_24 : bit_vector(255 downto 0) := X"7D7A7673706D6A6663605D5A5653504D4A4643403D3A3633302D2A2623201D1A";
constant INIT_H_HUM_25 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_HUM_25 : bit_vector(255 downto 0) := X"E3E0DDDAD6D3D0CDCAC6C3C0BDBAB6B3B0ADAAA6A3A09D9A9693908D8A868380";
constant INIT_H_HUM_26 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060505050505050505";
constant INIT_L_HUM_26 : bit_vector(255 downto 0) := X"4A4643403D3A3633302D2A2623201D1A1613100D0A060300FDFAF6F3F0EDEAE6";
constant INIT_H_HUM_27 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_HUM_27 : bit_vector(255 downto 0) := X"B0ADAAA6A3A09D9A9693908D8A8683807D7A7673706D6A6663605D5A5653504D";
constant INIT_H_HUM_28 : bit_vector(255 downto 0) := X"0707070707070707060606060606060606060606060606060606060606060606";
constant INIT_L_HUM_28 : bit_vector(255 downto 0) := X"1613100D09060300FDF9F6F3F0EDE9E6E3E0DDD9D6D3D0CDC9C6C3C0BDBAB6B3";
constant INIT_H_HUM_29 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_HUM_29 : bit_vector(255 downto 0) := X"7D797673706D696663605D595653504D494643403D393633302D292623201D19";
constant INIT_H_HUM_2A : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_HUM_2A : bit_vector(255 downto 0) := X"E3E0DDD9D6D3D0CDC9C6C3C0BDB9B6B3B0ADA9A6A3A09D999693908D89868380";
constant INIT_H_HUM_2B : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080707070707070707";
constant INIT_L_HUM_2B : bit_vector(255 downto 0) := X"494643403D393633302D292623201D191613100D09060300FDF9F6F3F0EDE9E6";
constant INIT_H_HUM_2C : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_HUM_2C : bit_vector(255 downto 0) := X"B0ADA9A6A3A09D999693908D898683807D797673706D696663605D595653504D";
constant INIT_H_HUM_2D : bit_vector(255 downto 0) := X"0909090909090909080808080808080808080808080808080808080808080808";
constant INIT_L_HUM_2D : bit_vector(255 downto 0) := X"1613100D09060300FDF9F6F3F0EDE9E6E3E0DDD9D6D3D0CDC9C6C3C0BDB9B6B3";
constant INIT_H_HUM_2E : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_HUM_2E : bit_vector(255 downto 0) := X"7D797673706D696663605D595653504D494643403D393633302D292623201D19";
constant INIT_H_HUM_2F : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_HUM_2F : bit_vector(255 downto 0) := X"E3E0DDD9D6D3D0CDC9C6C3C0BDB9B6B3B0ADA9A6A3A09D999693908D89868380";
constant INIT_H_HUM_30 : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0909090909090909";
constant INIT_L_HUM_30 : bit_vector(255 downto 0) := X"494643403D393633302D292623201D191613100D09060300FDF9F6F3F0EDE9E6";
constant INIT_H_HUM_31 : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_HUM_31 : bit_vector(255 downto 0) := X"B0ADA9A6A3A09D999693908D898683807D797673706D696663605D595653504D";
constant INIT_H_HUM_32 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_HUM_32 : bit_vector(255 downto 0) := X"1613100D09060300FDF9F6F3F0EDE9E6E3E0DDD9D6D3D0CDC9C6C3C0BDB9B6B3";
constant INIT_H_HUM_33 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_HUM_33 : bit_vector(255 downto 0) := X"7D797673706D696663605D595653504D494643403D393633302D292623201D19";
constant INIT_H_HUM_34 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_HUM_34 : bit_vector(255 downto 0) := X"E3E0DDD9D6D3D0CDC9C6C3C0BDB9B6B3B0ADA9A6A3A09D999693908D89868380";
constant INIT_H_HUM_35 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B0B";
constant INIT_L_HUM_35 : bit_vector(255 downto 0) := X"494643403D393633302D292623201D191613100D09060300FDF9F6F3F0EDE9E6";
constant INIT_H_HUM_36 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_HUM_36 : bit_vector(255 downto 0) := X"B0ADA9A6A3A09D999693908D898683807D797673706D696663605D595653504D";
constant INIT_H_HUM_37 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_HUM_37 : bit_vector(255 downto 0) := X"1613100D09060300FDF9F6F3F0EDE9E6E3E0DDD9D6D3D0CDC9C6C3C0BDB9B6B3";
constant INIT_H_HUM_38 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_HUM_38 : bit_vector(255 downto 0) := X"7D797673706D696663605D595653504D494643403D393633302D292623201D19";
constant INIT_H_HUM_39 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_HUM_39 : bit_vector(255 downto 0) := X"E3E0DDD9D6D3D0CDC9C6C3C0BDB9B6B3B0ADA9A6A3A09D999693908D89868380";
constant INIT_H_HUM_3A : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0D0D0D0D0D0D0D0D";
constant INIT_L_HUM_3A : bit_vector(255 downto 0) := X"494643403D393633302D292623201D191613100D09060300FDF9F6F3F0EDE9E6";
constant INIT_H_HUM_3B : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_HUM_3B : bit_vector(255 downto 0) := X"B0ADA9A6A3A09D999693908D898683807D797673706D696663605D595653504D";
constant INIT_H_HUM_3C : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_HUM_3C : bit_vector(255 downto 0) := X"1613100C09060300FCF9F6F3F0ECE9E6E3E0DCD9D6D3D0CCC9C6C3C0BDB9B6B3";
constant INIT_H_HUM_3D : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_HUM_3D : bit_vector(255 downto 0) := X"7C797673706C696663605C595653504C494643403C393633302C292623201C19";
constant INIT_H_HUM_3E : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_HUM_3E : bit_vector(255 downto 0) := X"E3E0DCD9D6D3D0CCC9C6C3C0BCB9B6B3B0ACA9A6A3A09C999693908C89868380";
constant INIT_H_HUM_3F : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010100F0F0F0F0F0F0F0F";
constant INIT_L_HUM_3F : bit_vector(255 downto 0) := X"494643403C393633302C292623201C191613100C09060300FCF9F6F3F0ECE9E6";
constant INIT_H_HUM_40 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_HUM_40 : bit_vector(255 downto 0) := X"B0ACA9A6A3A09C999693908C898683807C797673706C696663605C595653504C";
constant INIT_H_HUM_41 : bit_vector(255 downto 0) := X"1111111111111111101010101010101010101010101010101010101010101010";
constant INIT_L_HUM_41 : bit_vector(255 downto 0) := X"1613100C09060300FCF9F6F3F0ECE9E6E3E0DCD9D6D3D0CCC9C6C3C0BCB9B6B3";
constant INIT_H_HUM_42 : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_HUM_42 : bit_vector(255 downto 0) := X"7C797673706C696663605C595653504C494643403C393633302C292623201C19";
constant INIT_H_HUM_43 : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_HUM_43 : bit_vector(255 downto 0) := X"E3E0DCD9D6D3D0CCC9C6C3C0BCB9B6B3B0ACA9A6A3A09C999693908C89868380";
constant INIT_H_HUM_44 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121111111111111111";
constant INIT_L_HUM_44 : bit_vector(255 downto 0) := X"494643403C393633302C292623201C191613100C09060300FCF9F6F3F0ECE9E6";
constant INIT_H_HUM_45 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_HUM_45 : bit_vector(255 downto 0) := X"B0ACA9A6A3A09C999693908C898683807C797673706C696663605C595653504C";
constant INIT_H_HUM_46 : bit_vector(255 downto 0) := X"1313131313131313121212121212121212121212121212121212121212121212";
constant INIT_L_HUM_46 : bit_vector(255 downto 0) := X"1613100C09060300FCF9F6F3F0ECE9E6E3E0DCD9D6D3D0CCC9C6C3C0BCB9B6B3";
constant INIT_H_HUM_47 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_HUM_47 : bit_vector(255 downto 0) := X"7C797673706C696663605C595653504C494643403C393633302C292623201C19";
constant INIT_H_HUM_48 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_HUM_48 : bit_vector(255 downto 0) := X"E3E0DCD9D6D3D0CCC9C6C3C0BCB9B6B3B0ACA9A6A3A09C999693908C89868380";
constant INIT_H_HUM_49 : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141313131313131313";
constant INIT_L_HUM_49 : bit_vector(255 downto 0) := X"494643403C393633302C292623201C191613100C09060300FCF9F6F3F0ECE9E6";
constant INIT_H_HUM_4A : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_HUM_4A : bit_vector(255 downto 0) := X"B0ACA9A6A3A09C999693908C898683807C797673706C696663605C595653504C";
constant INIT_H_HUM_4B : bit_vector(255 downto 0) := X"1515151515151515141414141414141414141414141414141414141414141414";
constant INIT_L_HUM_4B : bit_vector(255 downto 0) := X"1613100C09060300FCF9F6F3F0ECE9E6E3E0DCD9D6D3D0CCC9C6C3C0BCB9B6B3";
constant INIT_H_HUM_4C : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_HUM_4C : bit_vector(255 downto 0) := X"7C797673706C696663605C595653504C494643403C393633302C292623201C19";
constant INIT_H_HUM_4D : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_HUM_4D : bit_vector(255 downto 0) := X"E3E0DCD9D6D3D0CCC9C6C3C0BCB9B6B3B0ACA9A6A3A09C999693908C89868380";
constant INIT_H_HUM_4E : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161515151515151515";
constant INIT_L_HUM_4E : bit_vector(255 downto 0) := X"494643403C393633302C292623201C191613100C09060300FCF9F6F3F0ECE9E6";
constant INIT_H_HUM_4F : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161616161616";
constant INIT_L_HUM_4F : bit_vector(255 downto 0) := X"B0ACA9A6A3A09C999693908C898683807C797673706C696663605C595653504C";
constant INIT_H_HUM_50 : bit_vector(255 downto 0) := X"1717171717171716161616161616161616161616161616161616161616161616";
constant INIT_L_HUM_50 : bit_vector(255 downto 0) := X"16130F0C090603FFFCF9F6F3EFECE9E6E3DFDCD9D6D3CFCCC9C6C3C0BCB9B6B3";
constant INIT_H_HUM_51 : bit_vector(255 downto 0) := X"1717171717171717171717171717171717171717171717171717171717171717";
constant INIT_L_HUM_51 : bit_vector(255 downto 0) := X"7C7976736F6C6966635F5C5956534F4C4946433F3C3936332F2C2926231F1C19";
constant INIT_H_HUM_52 : bit_vector(255 downto 0) := X"1717171717171717171717171717171717171717171717171717171717171717";
constant INIT_L_HUM_52 : bit_vector(255 downto 0) := X"E3DFDCD9D6D3CFCCC9C6C3BFBCB9B6B3AFACA9A6A39F9C9996938F8C8986837F";
constant INIT_H_HUM_53 : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818171717171717171717";
constant INIT_L_HUM_53 : bit_vector(255 downto 0) := X"4946433F3C3936332F2C2926231F1C1916130F0C090603FFFCF9F6F3EFECE9E6";
constant INIT_H_HUM_54 : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_HUM_54 : bit_vector(255 downto 0) := X"AFACA9A6A39F9C9996938F8C8986837F7C7976736F6C6966635F5C5956534F4C";
constant INIT_H_HUM_55 : bit_vector(255 downto 0) := X"1919191919191918181818181818181818181818181818181818181818181818";
constant INIT_L_HUM_55 : bit_vector(255 downto 0) := X"16130F0C090603FFFCF9F6F3EFECE9E6E3DFDCD9D6D3CFCCC9C6C3BFBCB9B6B3";
constant INIT_H_HUM_56 : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_HUM_56 : bit_vector(255 downto 0) := X"7C7976736F6C6966635F5C5956534F4C4946433F3C3936332F2C2926231F1C19";
constant INIT_H_HUM_57 : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_HUM_57 : bit_vector(255 downto 0) := X"E3DFDCD9D6D3CFCCC9C6C3BFBCB9B6B3AFACA9A6A39F9C9996938F8C8986837F";
constant INIT_H_HUM_58 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A191919191919191919";
constant INIT_L_HUM_58 : bit_vector(255 downto 0) := X"4946433F3C3936332F2C2926231F1C1916130F0C090603FFFCF9F6F3EFECE9E6";
constant INIT_H_HUM_59 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_HUM_59 : bit_vector(255 downto 0) := X"AFACA9A6A39F9C9996938F8C8986837F7C7976736F6C6966635F5C5956534F4C";
constant INIT_H_HUM_5A : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_HUM_5A : bit_vector(255 downto 0) := X"16130F0C090603FFFCF9F6F3EFECE9E6E3DFDCD9D6D3CFCCC9C6C3BFBCB9B6B3";
constant INIT_H_HUM_5B : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_HUM_5B : bit_vector(255 downto 0) := X"7C7976736F6C6966635F5C5956534F4C4946433F3C3936332F2C2926231F1C19";
constant INIT_H_HUM_5C : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_HUM_5C : bit_vector(255 downto 0) := X"E3DFDCD9D6D3CFCCC9C6C3BFBCB9B6B3AFACA9A6A39F9C9996938F8C8986837F";
constant INIT_H_HUM_5D : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1B1B1B1B1B1B1B1B1B";
constant INIT_L_HUM_5D : bit_vector(255 downto 0) := X"4946433F3C3936332F2C2926231F1C1916130F0C090603FFFCF9F6F3EFECE9E6";
constant INIT_H_HUM_5E : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_HUM_5E : bit_vector(255 downto 0) := X"AFACA9A6A39F9C9996938F8C8986837F7C7976736F6C6966635F5C5956534F4C";
constant INIT_H_HUM_5F : bit_vector(255 downto 0) := X"1D1D1D1D1D1D1D1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_HUM_5F : bit_vector(255 downto 0) := X"16130F0C090603FFFCF9F6F3EFECE9E6E3DFDCD9D6D3CFCCC9C6C3BFBCB9B6B3";
constant INIT_H_HUM_60 : bit_vector(255 downto 0) := X"1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D";
constant INIT_L_HUM_60 : bit_vector(255 downto 0) := X"7C7976736F6C6966635F5C5956534F4C4946433F3C3936332F2C2926231F1C19";
constant INIT_H_HUM_61 : bit_vector(255 downto 0) := X"1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D";
constant INIT_L_HUM_61 : bit_vector(255 downto 0) := X"E3DFDCD9D6D3CFCCC9C6C3BFBCB9B6B3AFACA9A6A39F9C9996938F8C8986837F";
constant INIT_H_HUM_62 : bit_vector(255 downto 0) := X"1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1D1D1D1D1D1D1D1D1D";
constant INIT_L_HUM_62 : bit_vector(255 downto 0) := X"4946433F3C3936332F2C2926231F1C1916130F0C090603FFFCF9F6F3EFECE9E6";
constant INIT_H_HUM_63 : bit_vector(255 downto 0) := X"1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E";
constant INIT_L_HUM_63 : bit_vector(255 downto 0) := X"AFACA9A6A39F9C9996938F8C8986837F7C7976736F6C6966635F5C5956534F4C";
constant INIT_H_HUM_64 : bit_vector(255 downto 0) := X"1F1F1F1F1F1F1F1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E";
constant INIT_L_HUM_64 : bit_vector(255 downto 0) := X"16120F0C090602FFFCF9F6F2EFECE9E6E2DFDCD9D6D2CFCCC9C6C3BFBCB9B6B3";
constant INIT_H_HUM_65 : bit_vector(255 downto 0) := X"1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F";
constant INIT_L_HUM_65 : bit_vector(255 downto 0) := X"7C7976726F6C6966625F5C5956524F4C4946423F3C3936322F2C2926221F1C19";
constant INIT_H_HUM_66 : bit_vector(255 downto 0) := X"1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F";
constant INIT_L_HUM_66 : bit_vector(255 downto 0) := X"E2DFDCD9D6D2CFCCC9C6C2BFBCB9B6B2AFACA9A6A29F9C9996928F8C8986827F";
constant INIT_H_HUM_67 : bit_vector(255 downto 0) := X"20202020202020202020202020202020202020202020201F1F1F1F1F1F1F1F1F";
constant INIT_L_HUM_67 : bit_vector(255 downto 0) := X"4946423F3C3936322F2C2926221F1C1916120F0C090602FFFCF9F6F2EFECE9E6";
constant INIT_H_HUM_68 : bit_vector(255 downto 0) := X"2020202020202020202020202020202020202020202020202020202020202020";
constant INIT_L_HUM_68 : bit_vector(255 downto 0) := X"AFACA9A6A29F9C9996928F8C8986827F7C7976726F6C6966625F5C5956524F4C";
constant INIT_H_HUM_69 : bit_vector(255 downto 0) := X"2121212121212120202020202020202020202020202020202020202020202020";
constant INIT_L_HUM_69 : bit_vector(255 downto 0) := X"16120F0C090602FFFCF9F6F2EFECE9E6E2DFDCD9D6D2CFCCC9C6C2BFBCB9B6B2";
constant INIT_H_HUM_6A : bit_vector(255 downto 0) := X"2121212121212121212121212121212121212121212121212121212121212121";
constant INIT_L_HUM_6A : bit_vector(255 downto 0) := X"7C7976726F6C6966625F5C5956524F4C4946423F3C3936322F2C2926221F1C19";
constant INIT_H_HUM_6B : bit_vector(255 downto 0) := X"2121212121212121212121212121212121212121212121212121212121212121";
constant INIT_L_HUM_6B : bit_vector(255 downto 0) := X"E2DFDCD9D6D2CFCCC9C6C2BFBCB9B6B2AFACA9A6A29F9C9996928F8C8986827F";
constant INIT_H_HUM_6C : bit_vector(255 downto 0) := X"2222222222222222222222222222222222222222222222212121212121212121";
constant INIT_L_HUM_6C : bit_vector(255 downto 0) := X"4946423F3C3936322F2C2926221F1C1916120F0C090602FFFCF9F6F2EFECE9E6";
constant INIT_H_HUM_6D : bit_vector(255 downto 0) := X"2222222222222222222222222222222222222222222222222222222222222222";
constant INIT_L_HUM_6D : bit_vector(255 downto 0) := X"AFACA9A6A29F9C9996928F8C8986827F7C7976726F6C6966625F5C5956524F4C";
constant INIT_H_HUM_6E : bit_vector(255 downto 0) := X"2323232323232322222222222222222222222222222222222222222222222222";
constant INIT_L_HUM_6E : bit_vector(255 downto 0) := X"16120F0C090602FFFCF9F6F2EFECE9E6E2DFDCD9D6D2CFCCC9C6C2BFBCB9B6B2";
constant INIT_H_HUM_6F : bit_vector(255 downto 0) := X"2323232323232323232323232323232323232323232323232323232323232323";
constant INIT_L_HUM_6F : bit_vector(255 downto 0) := X"7C7976726F6C6966625F5C5956524F4C4946423F3C3936322F2C2926221F1C19";
constant INIT_H_HUM_70 : bit_vector(255 downto 0) := X"2323232323232323232323232323232323232323232323232323232323232323";
constant INIT_L_HUM_70 : bit_vector(255 downto 0) := X"E2DFDCD9D6D2CFCCC9C6C2BFBCB9B6B2AFACA9A6A29F9C9996928F8C8986827F";
constant INIT_H_HUM_71 : bit_vector(255 downto 0) := X"2424242424242424242424242424242424242424242424232323232323232323";
constant INIT_L_HUM_71 : bit_vector(255 downto 0) := X"4946423F3C3936322F2C2926221F1C1916120F0C090602FFFCF9F6F2EFECE9E6";
constant INIT_H_HUM_72 : bit_vector(255 downto 0) := X"2424242424242424242424242424242424242424242424242424242424242424";
constant INIT_L_HUM_72 : bit_vector(255 downto 0) := X"AFACA9A6A29F9C9996928F8C8986827F7C7976726F6C6966625F5C5956524F4C";
constant INIT_H_HUM_73 : bit_vector(255 downto 0) := X"2525252525252524242424242424242424242424242424242424242424242424";
constant INIT_L_HUM_73 : bit_vector(255 downto 0) := X"16120F0C090602FFFCF9F6F2EFECE9E6E2DFDCD9D6D2CFCCC9C6C2BFBCB9B6B2";
constant INIT_H_HUM_74 : bit_vector(255 downto 0) := X"2525252525252525252525252525252525252525252525252525252525252525";
constant INIT_L_HUM_74 : bit_vector(255 downto 0) := X"7C7976726F6C6966625F5C5956524F4C4946423F3C3936322F2C2926221F1C19";
constant INIT_H_HUM_75 : bit_vector(255 downto 0) := X"2525252525252525252525252525252525252525252525252525252525252525";
constant INIT_L_HUM_75 : bit_vector(255 downto 0) := X"E2DFDCD9D6D2CFCCC9C6C2BFBCB9B6B2AFACA9A6A29F9C9996928F8C8986827F";
constant INIT_H_HUM_76 : bit_vector(255 downto 0) := X"2626262626262626262626262626262626262626262626252525252525252525";
constant INIT_L_HUM_76 : bit_vector(255 downto 0) := X"4946423F3C3936322F2C2926221F1C1916120F0C090602FFFCF9F6F2EFECE9E6";
constant INIT_H_HUM_77 : bit_vector(255 downto 0) := X"2626262626262626262626262626262626262626262626262626262626262626";
constant INIT_L_HUM_77 : bit_vector(255 downto 0) := X"AFACA9A6A29F9C9996928F8C8986827F7C7976726F6C6966625F5C5956524F4C";
constant INIT_H_HUM_78 : bit_vector(255 downto 0) := X"2727272727272726262626262626262626262626262626262626262626262626";
constant INIT_L_HUM_78 : bit_vector(255 downto 0) := X"15120F0C090502FFFCF9F5F2EFECE9E5E2DFDCD9D5D2CFCCC9C6C2BFBCB9B6B2";
constant INIT_H_HUM_79 : bit_vector(255 downto 0) := X"2727272727272727272727272727272727272727272727272727272727272727";
constant INIT_L_HUM_79 : bit_vector(255 downto 0) := X"7C7975726F6C6965625F5C5955524F4C4945423F3C3935322F2C2925221F1C19";
constant INIT_H_HUM_7A : bit_vector(255 downto 0) := X"2727272727272727272727272727272727272727272727272727272727272727";
constant INIT_L_HUM_7A : bit_vector(255 downto 0) := X"E2DFDCD9D5D2CFCCC9C5C2BFBCB9B5B2AFACA9A5A29F9C9995928F8C8985827F";
constant INIT_H_HUM_7B : bit_vector(255 downto 0) := X"2828282828282828282828282828282828282828282828272727272727272727";
constant INIT_L_HUM_7B : bit_vector(255 downto 0) := X"4945423F3C3935322F2C2925221F1C1915120F0C090502FFFCF9F5F2EFECE9E5";
constant INIT_H_HUM_7C : bit_vector(255 downto 0) := X"2828282828282828282828282828282828282828282828282828282828282828";
constant INIT_L_HUM_7C : bit_vector(255 downto 0) := X"AFACA9A5A29F9C9995928F8C8985827F7C7975726F6C6965625F5C5955524F4C";
constant INIT_H_HUM_7D : bit_vector(255 downto 0) := X"2929292929292928282828282828282828282828282828282828282828282828";
constant INIT_L_HUM_7D : bit_vector(255 downto 0) := X"15120F0C090502FFFCF9F5F2EFECE9E5E2DFDCD9D5D2CFCCC9C5C2BFBCB9B5B2";
constant INIT_H_HUM_7E : bit_vector(255 downto 0) := X"2929292929292929292929292929292929292929292929292929292929292929";
constant INIT_L_HUM_7E : bit_vector(255 downto 0) := X"7C7975726F6C6965625F5C5955524F4C4945423F3C3935322F2C2925221F1C19";
constant INIT_H_HUM_7F : bit_vector(255 downto 0) := X"2929292929292929292929292929292929292929292929292929292929292929";
constant INIT_L_HUM_7F : bit_vector(255 downto 0) := X"E2DFDCD9D5D2CFCCC9C5C2BFBCB9B5B2AFACA9A5A29F9C9995928F8C8985827F";
constant INIT_H_IANA_00 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IANA_00 : bit_vector(255 downto 0) := X"504D4B484643403E3B393633312E2C292624211F1C191714120F0C0A07050200";
constant INIT_H_IANA_01 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IANA_01 : bit_vector(255 downto 0) := X"A3A19E9B999694918E8C898784817F7C7A7774726F6D6A676562605D5A585553";
constant INIT_H_IANA_02 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IANA_02 : bit_vector(255 downto 0) := X"F6F4F1EFECE9E7E4E2DFDCDAD7D5D2CFCDCAC8C5C2C0BDBBB8B5B3B0AEABA8A6";
constant INIT_H_IANA_03 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101000000";
constant INIT_L_IANA_03 : bit_vector(255 downto 0) := X"494744423F3C3A3735322F2D2A282522201D1B181513100E0B08060301FEFBF9";
constant INIT_H_IANA_04 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IANA_04 : bit_vector(255 downto 0) := X"9D9A979592908D8A888583807D7B787673706E6B696663615E5C595654514F4C";
constant INIT_H_IANA_05 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IANA_05 : bit_vector(255 downto 0) := X"F0EDEAE8E5E3E0DEDBD8D6D3D1CECBC9C6C4C1BEBCB9B7B4B1AFACAAA7A4A29F";
constant INIT_H_IANA_06 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202010101010101";
constant INIT_L_IANA_06 : bit_vector(255 downto 0) := X"43403E3B383633312E2B292624211E1C191714110F0C0A070402FFFDFAF7F5F2";
constant INIT_H_IANA_07 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IANA_07 : bit_vector(255 downto 0) := X"9693918E8C898684817F7C797774726F6C6A6765625F5D5A585552504D4B4845";
constant INIT_H_IANA_08 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IANA_08 : bit_vector(255 downto 0) := X"E9E6E4E1DFDCDAD7D4D2CFCDCAC7C5C2C0BDBAB8B5B3B0ADABA8A6A3A09E9B99";
constant INIT_H_IANA_09 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030202020202020202";
constant INIT_L_IANA_09 : bit_vector(255 downto 0) := X"3C3A3734322F2D2A272522201D1A181513100D0B08060300FEFBF9F6F3F1EEEC";
constant INIT_H_IANA_0A : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IANA_0A : bit_vector(255 downto 0) := X"8F8D8A888582807D7B787573706E6B686663615E5B595654514E4C494744413F";
constant INIT_H_IANA_0B : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IANA_0B : bit_vector(255 downto 0) := X"E2E0DDDBD8D5D3D0CECBC9C6C3C1BEBCB9B6B4B1AFACA9A7A4A29F9C9A979592";
constant INIT_H_IANA_0C : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040303030303030303030303";
constant INIT_L_IANA_0C : bit_vector(255 downto 0) := X"3633302E2B292623211E1C191614110F0C09070402FFFCFAF7F5F2EFEDEAE8E5";
constant INIT_H_IANA_0D : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IANA_0D : bit_vector(255 downto 0) := X"898684817E7C797774716F6C6A6764625F5D5A575552504D4A484543403D3B38";
constant INIT_H_IANA_0E : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IANA_0E : bit_vector(255 downto 0) := X"DCD9D7D4D1CFCCCAC7C5C2BFBDBAB8B5B2B0ADABA8A5A3A09E9B989693918E8B";
constant INIT_H_IANA_0F : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050504040404040404040404040404";
constant INIT_L_IANA_0F : bit_vector(255 downto 0) := X"2F2C2A2725221F1D1A181512100D0B08050300FEFBF8F6F3F1EEEBE9E6E4E1DE";
constant INIT_H_IANA_10 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IANA_10 : bit_vector(255 downto 0) := X"82807D7A787573706D6B686663605E5B595653514E4C494644413F3C39373432";
constant INIT_H_IANA_11 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IANA_11 : bit_vector(255 downto 0) := X"D5D3D0CDCBC8C6C3C0BEBBB9B6B4B1AEACA9A7A4A19F9C9A9794928F8D8A8785";
constant INIT_H_IANA_12 : bit_vector(255 downto 0) := X"0606060606060606060606060606060605050505050505050505050505050505";
constant INIT_L_IANA_12 : bit_vector(255 downto 0) := X"282623211E1B191614110E0C09070401FFFCFAF7F4F2EFEDEAE7E5E2E0DDDAD8";
constant INIT_H_IANA_13 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IANA_13 : bit_vector(255 downto 0) := X"7C797674716F6C696764625F5C5A5755524F4D4A484542403D3B383533302E2B";
constant INIT_H_IANA_14 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IANA_14 : bit_vector(255 downto 0) := X"CFCCC9C7C4C2BFBCBAB7B5B2AFADAAA8A5A3A09D9B989693908E8B898683817E";
constant INIT_H_IANA_15 : bit_vector(255 downto 0) := X"0707070707070707070707070707060606060606060606060606060606060606";
constant INIT_L_IANA_15 : bit_vector(255 downto 0) := X"221F1D1A171512100D0A08050300FDFBF8F6F3F0EEEBE9E6E3E1DEDCD9D6D4D1";
constant INIT_H_IANA_16 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IANA_16 : bit_vector(255 downto 0) := X"7572706D6B686563605E5B585653514E4B494644413E3C393734312F2C2A2724";
constant INIT_H_IANA_17 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IANA_17 : bit_vector(255 downto 0) := X"C8C5C3C0BEBBB8B6B3B1AEABA9A6A4A19F9C999794928F8C8A8785827F7D7A78";
constant INIT_H_IANA_18 : bit_vector(255 downto 0) := X"0808080808080808080808070707070707070707070707070707070707070707";
constant INIT_L_IANA_18 : bit_vector(255 downto 0) := X"1B191613110E0C09060401FFFCF9F7F4F2EFECEAE7E5E2DFDDDAD8D5D2D0CDCB";
constant INIT_H_IANA_19 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IANA_19 : bit_vector(255 downto 0) := X"6E6C696764615F5C5A5754524F4D4A474542403D3A383533302D2B282623201E";
constant INIT_H_IANA_1A : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IANA_1A : bit_vector(255 downto 0) := X"C1BFBCBAB7B4B2AFADAAA7A5A2A09D9A989593908E8B888683817E7B79767471";
constant INIT_H_IANA_1B : bit_vector(255 downto 0) := X"0909090909090909090808080808080808080808080808080808080808080808";
constant INIT_L_IANA_1B : bit_vector(255 downto 0) := X"15120F0D0A08050200FDFBF8F5F3F0EEEBE8E6E3E1DEDBD9D6D4D1CECCC9C7C4";
constant INIT_H_IANA_1C : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IANA_1C : bit_vector(255 downto 0) := X"686563605D5B585653504E4B494643413E3C393634312F2C292724221F1C1A17";
constant INIT_H_IANA_1D : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IANA_1D : bit_vector(255 downto 0) := X"BBB8B6B3B0AEABA9A6A3A19E9C999694918F8C8A8784827F7D7A777572706D6A";
constant INIT_H_IANA_1E : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0909090909090909090909090909090909090909090909090909";
constant INIT_L_IANA_1E : bit_vector(255 downto 0) := X"0E0B09060401FEFCF9F7F4F1EFECEAE7E4E2DFDDDAD7D5D2D0CDCAC8C5C3C0BD";
constant INIT_H_IANA_1F : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_IANA_1F : bit_vector(255 downto 0) := X"615F5C595754524F4C4A4745423F3D3A383532302D2B282523201E1B18161311";
constant INIT_H_IANA_20 : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_IANA_20 : bit_vector(255 downto 0) := X"B4B2AFACAAA7A5A29F9D9A989592908D8B888583807E7B797673716E6C696664";
constant INIT_H_IANA_21 : bit_vector(255 downto 0) := X"0B0B0B0B0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_IANA_21 : bit_vector(255 downto 0) := X"07050200FDFAF8F5F3F0EDEBE8E6E3E0DEDBD9D6D3D1CECCC9C6C4C1BFBCB9B7";
constant INIT_H_IANA_22 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_IANA_22 : bit_vector(255 downto 0) := X"5B585553504E4B484643413E3B393634312E2C292724211F1C1A1714120F0D0A";
constant INIT_H_IANA_23 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_IANA_23 : bit_vector(255 downto 0) := X"AEABA8A6A3A19E9B999694918E8C898784817F7C7A7775726F6D6A686562605D";
constant INIT_H_IANA_24 : bit_vector(255 downto 0) := X"0C0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_IANA_24 : bit_vector(255 downto 0) := X"01FEFCF9F6F4F1EFECE9E7E4E2DFDCDAD7D5D2CFCDCAC8C5C2C0BDBBB8B5B3B0";
constant INIT_H_IANA_25 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_IANA_25 : bit_vector(255 downto 0) := X"54514F4C4A4744423F3D3A373532302D2A282523201D1B181613100E0B090603";
constant INIT_H_IANA_26 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_IANA_26 : bit_vector(255 downto 0) := X"A7A4A29F9D9A979592908D8A888583807D7B787673706E6B696664615E5C5957";
constant INIT_H_IANA_27 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_IANA_27 : bit_vector(255 downto 0) := X"FAF8F5F2F0EDEBE8E5E3E0DEDBD8D6D3D1CECBC9C6C4C1BEBCB9B7B4B1AFACAA";
constant INIT_H_IANA_28 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0C0C";
constant INIT_L_IANA_28 : bit_vector(255 downto 0) := X"4D4B484643403E3B393633312E2C292624211F1C191714120F0C0A070502FFFD";
constant INIT_H_IANA_29 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_IANA_29 : bit_vector(255 downto 0) := X"A09E9B999693918E8C898684817F7C797774726F6C6A6765625F5D5A58555350";
constant INIT_H_IANA_2A : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_IANA_2A : bit_vector(255 downto 0) := X"F4F1EEECE9E7E4E1DFDCDAD7D4D2CFCDCAC7C5C2C0BDBAB8B5B3B0ADABA8A6A3";
constant INIT_H_IANA_2B : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0D0D0D0D";
constant INIT_L_IANA_2B : bit_vector(255 downto 0) := X"4744423F3C3A3735322F2D2A282522201D1B181513100E0B08060301FEFBF9F6";
constant INIT_H_IANA_2C : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_IANA_2C : bit_vector(255 downto 0) := X"9A9795928F8D8A888582807D7B787573706E6B686663615E5B595654514F4C49";
constant INIT_H_IANA_2D : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_IANA_2D : bit_vector(255 downto 0) := X"EDEAE8E5E3E0DDDBD8D6D3D0CECBC9C6C3C1BEBCB9B6B4B1AFACA9A7A4A29F9C";
constant INIT_H_IANA_2E : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0E0E0E0E0E0E0E";
constant INIT_L_IANA_2E : bit_vector(255 downto 0) := X"403E3B383633312E2B292624211E1C191714110F0C0A070402FFFDFAF7F5F2F0";
constant INIT_H_IANA_2F : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_IANA_2F : bit_vector(255 downto 0) := X"93918E8B898684817E7C797774716F6C6A6764625F5D5A575552504D4A484543";
constant INIT_H_IANA_30 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_IANA_30 : bit_vector(255 downto 0) := X"E6E4E1DFDCD9D7D4D2CFCCCAC7C5C2BFBDBAB8B5B2B0ADABA8A5A3A09E9B9896";
constant INIT_H_IANA_31 : bit_vector(255 downto 0) := X"10101010101010101010101010101010101010101010100F0F0F0F0F0F0F0F0F";
constant INIT_L_IANA_31 : bit_vector(255 downto 0) := X"3A3734322F2D2A272522201D1A181513100D0B08060300FEFBF9F6F3F1EEECE9";
constant INIT_H_IANA_32 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_IANA_32 : bit_vector(255 downto 0) := X"8D8A878582807D7A787573706D6B686663605E5B595653514E4C494644413F3C";
constant INIT_H_IANA_33 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_IANA_33 : bit_vector(255 downto 0) := X"E0DDDBD8D5D3D0CECBC8C6C3C1BEBBB9B6B4B1AEACA9A7A4A19F9C9A9794928F";
constant INIT_H_IANA_34 : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111101010101010101010101010";
constant INIT_L_IANA_34 : bit_vector(255 downto 0) := X"33302E2B292623211E1C191614110F0C09070402FFFCFAF7F5F2EFEDEAE8E5E2";
constant INIT_H_IANA_35 : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_IANA_35 : bit_vector(255 downto 0) := X"8683817E7C797674716F6C696764625F5C5A5755524F4D4A484542403D3B3835";
constant INIT_H_IANA_36 : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_IANA_36 : bit_vector(255 downto 0) := X"D9D7D4D1CFCCCAC7C4C2BFBDBAB7B5B2B0ADAAA8A5A3A09D9B989693908E8B89";
constant INIT_H_IANA_37 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121111111111111111111111111111";
constant INIT_L_IANA_37 : bit_vector(255 downto 0) := X"2C2A2725221F1D1A181512100D0B08050300FEFBF8F6F3F1EEEBE9E6E4E1DEDC";
constant INIT_H_IANA_38 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_IANA_38 : bit_vector(255 downto 0) := X"7F7D7A787572706D6B686563605E5B585653514E4B494644413E3C393734312F";
constant INIT_H_IANA_39 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_IANA_39 : bit_vector(255 downto 0) := X"D3D0CDCBC8C6C3C0BEBBB9B6B3B1AEACA9A6A4A19F9C999794928F8C8A878582";
constant INIT_H_IANA_3A : bit_vector(255 downto 0) := X"1313131313131313131313131313131212121212121212121212121212121212";
constant INIT_L_IANA_3A : bit_vector(255 downto 0) := X"2623201E1B191614110E0C09070401FFFCFAF7F4F2EFEDEAE7E5E2E0DDDAD8D5";
constant INIT_H_IANA_3B : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_IANA_3B : bit_vector(255 downto 0) := X"797674716E6C696764615F5C5A5754524F4D4A474542403D3A383533302D2B28";
constant INIT_H_IANA_3C : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_IANA_3C : bit_vector(255 downto 0) := X"CCC9C7C4C2BFBCBAB7B5B2AFADAAA8A5A2A09D9B989593908E8B888683817E7B";
constant INIT_H_IANA_3D : bit_vector(255 downto 0) := X"1414141414141414141414141413131313131313131313131313131313131313";
constant INIT_L_IANA_3D : bit_vector(255 downto 0) := X"1F1C1A1715120F0D0A08050300FDFBF8F6F3F0EEEBE9E6E3E1DEDCD9D6D4D1CF";
constant INIT_H_IANA_3E : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_IANA_3E : bit_vector(255 downto 0) := X"72706D6A686563605D5B585653504E4B494643413E3C393634312F2C29272422";
constant INIT_H_IANA_3F : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_IANA_3F : bit_vector(255 downto 0) := X"C5C3C0BEBBB8B6B3B1AEABA9A6A4A19E9C999794918F8C8A8784827F7D7A7775";
constant INIT_H_IANA_40 : bit_vector(255 downto 0) := X"1515151515151515151514141414141414141414141414141414141414141414";
constant INIT_L_IANA_40 : bit_vector(255 downto 0) := X"181613110E0B09060401FFFCF9F7F4F2EFECEAE7E5E2DFDDDAD8D5D2D0CDCBC8";
constant INIT_H_IANA_41 : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_IANA_41 : bit_vector(255 downto 0) := X"6C696664615F5C595754524F4C4A4745423F3D3A383532302D2B282523201E1B";
constant INIT_H_IANA_42 : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_IANA_42 : bit_vector(255 downto 0) := X"BFBCBAB7B4B2AFADAAA7A5A2A09D9A989593908D8B888683807E7B797673716E";
constant INIT_H_IANA_43 : bit_vector(255 downto 0) := X"1616161616161616151515151515151515151515151515151515151515151515";
constant INIT_L_IANA_43 : bit_vector(255 downto 0) := X"120F0D0A07050200FDFAF8F5F3F0EEEBE8E6E3E1DEDBD9D6D4D1CECCC9C7C4C1";
constant INIT_H_IANA_44 : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161616161616";
constant INIT_L_IANA_44 : bit_vector(255 downto 0) := X"6562605D5B585553504E4B484643413E3B393634312E2C292724211F1C1A1714";
constant INIT_H_IANA_45 : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161616161616";
constant INIT_L_IANA_45 : bit_vector(255 downto 0) := X"B8B6B3B0AEABA9A6A3A19E9C999694918F8C898784827F7C7A7775726F6D6A68";
constant INIT_H_IANA_46 : bit_vector(255 downto 0) := X"1717171717161616161616161616161616161616161616161616161616161616";
constant INIT_L_IANA_46 : bit_vector(255 downto 0) := X"0B09060301FEFCF9F6F4F1EFECEAE7E4E2DFDDDAD7D5D2D0CDCAC8C5C3C0BDBB";
constant INIT_H_IANA_47 : bit_vector(255 downto 0) := X"1717171717171717171717171717171717171717171717171717171717171717";
constant INIT_L_IANA_47 : bit_vector(255 downto 0) := X"5E5C595754514F4C4A4744423F3D3A373532302D2A282523201D1B181613100E";
constant INIT_H_IANA_48 : bit_vector(255 downto 0) := X"1717171717171717171717171717171717171717171717171717171717171717";
constant INIT_L_IANA_48 : bit_vector(255 downto 0) := X"B2AFACAAA7A5A29F9D9A989592908D8B888583807E7B787673716E6B69666461";
constant INIT_H_IANA_49 : bit_vector(255 downto 0) := X"1818171717171717171717171717171717171717171717171717171717171717";
constant INIT_L_IANA_49 : bit_vector(255 downto 0) := X"0502FFFDFAF8F5F2F0EDEBE8E5E3E0DEDBD9D6D3D1CECCC9C6C4C1BFBCB9B7B4";
constant INIT_H_IANA_4A : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_IANA_4A : bit_vector(255 downto 0) := X"585553504D4B484643403E3B393633312E2C292624211F1C191714120F0C0A07";
constant INIT_H_IANA_4B : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_IANA_4B : bit_vector(255 downto 0) := X"ABA8A6A3A19E9B999694918E8C898784817F7C7A7774726F6D6A676562605D5A";
constant INIT_H_IANA_4C : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_IANA_4C : bit_vector(255 downto 0) := X"FEFBF9F6F4F1EEECE9E7E4E1DFDCDAD7D5D2CFCDCAC8C5C2C0BDBBB8B5B3B0AE";
constant INIT_H_IANA_4D : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_IANA_4D : bit_vector(255 downto 0) := X"514F4C494744423F3C3A3735322F2D2A282522201D1B181513100E0B08060301";
constant INIT_H_IANA_4E : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_IANA_4E : bit_vector(255 downto 0) := X"A4A29F9D9A979592908D8A888583807D7B787673706E6B696663615E5C595654";
constant INIT_H_IANA_4F : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_IANA_4F : bit_vector(255 downto 0) := X"F7F5F2F0EDEAE8E5E3E0DDDBD8D6D3D0CECBC9C6C4C1BEBCB9B7B4B1AFACAAA7";
constant INIT_H_IANA_50 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A191919";
constant INIT_L_IANA_50 : bit_vector(255 downto 0) := X"4B484543403E3B383633312E2B292624211E1C191714110F0C0A070402FFFDFA";
constant INIT_H_IANA_51 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_IANA_51 : bit_vector(255 downto 0) := X"9E9B999693918E8C898684817F7C797774726F6C6A6765625F5D5A585552504D";
constant INIT_H_IANA_52 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_IANA_52 : bit_vector(255 downto 0) := X"F1EEECE9E6E4E1DFDCD9D7D4D2CFCCCAC7C5C2BFBDBAB8B5B3B0ADABA8A6A3A0";
constant INIT_H_IANA_53 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1A1A1A1A1A";
constant INIT_L_IANA_53 : bit_vector(255 downto 0) := X"44413F3C3A3734322F2D2A272522201D1A181513100D0B08060300FEFBF9F6F3";
constant INIT_H_IANA_54 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_IANA_54 : bit_vector(255 downto 0) := X"9795928F8D8A888582807D7B787573706E6B686663615E5B595654514E4C4947";
constant INIT_H_IANA_55 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_IANA_55 : bit_vector(255 downto 0) := X"EAE8E5E2E0DDDBD8D5D3D0CECBC8C6C3C1BEBBB9B6B4B1AFACA9A7A4A29F9C9A";
constant INIT_H_IANA_56 : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1B1B1B1B1B1B1B1B";
constant INIT_L_IANA_56 : bit_vector(255 downto 0) := X"3D3B383633302E2B292623211E1C191614110F0C09070402FFFCFAF7F5F2EFED";
constant INIT_H_IANA_57 : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_IANA_57 : bit_vector(255 downto 0) := X"918E8B898684817E7C797774716F6C6A6764625F5D5A575552504D4A48454340";
constant INIT_H_IANA_58 : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_IANA_58 : bit_vector(255 downto 0) := X"E4E1DEDCD9D7D4D1CFCCCAC7C4C2BFBDBAB7B5B2B0ADAAA8A5A3A09E9B989693";
constant INIT_H_IANA_59 : bit_vector(255 downto 0) := X"1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_IANA_59 : bit_vector(255 downto 0) := X"3734322F2C2A2725221F1D1A181512100D0B08050300FEFBF8F6F3F1EEEBE9E6";
constant INIT_H_IANA_5A : bit_vector(255 downto 0) := X"1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D";
constant INIT_L_IANA_5A : bit_vector(255 downto 0) := X"8A878582807D7A787573706D6B686663605E5B595653514E4C494644413F3C39";
constant INIT_H_IANA_5B : bit_vector(255 downto 0) := X"1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D";
constant INIT_L_IANA_5B : bit_vector(255 downto 0) := X"DDDAD8D5D3D0CDCBC8C6C3C0BEBBB9B6B3B1AEACA9A6A4A19F9C9A9794928F8D";
constant INIT_H_IANA_5C : bit_vector(255 downto 0) := X"1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1D1D1D1D1D1D1D1D1D1D1D1D1D";
constant INIT_L_IANA_5C : bit_vector(255 downto 0) := X"302E2B282623211E1B191614110E0C09070401FFFCFAF7F4F2EFEDEAE7E5E2E0";
constant INIT_H_IANA_5D : bit_vector(255 downto 0) := X"1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E";
constant INIT_L_IANA_5D : bit_vector(255 downto 0) := X"83817E7C797674716F6C696764625F5C5A5755524F4D4A484542403D3B383533";
constant INIT_H_IANA_5E : bit_vector(255 downto 0) := X"1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E";
constant INIT_L_IANA_5E : bit_vector(255 downto 0) := X"D6D4D1CFCCC9C7C4C2BFBCBAB7B5B2AFADAAA8A5A2A09D9B989593908E8B8986";
constant INIT_H_IANA_5F : bit_vector(255 downto 0) := X"1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E";
constant INIT_L_IANA_5F : bit_vector(255 downto 0) := X"2A2724221F1D1A171512100D0A08050300FDFBF8F6F3F0EEEBE9E6E3E1DEDCD9";
constant INIT_H_IANA_60 : bit_vector(255 downto 0) := X"1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F";
constant INIT_L_IANA_60 : bit_vector(255 downto 0) := X"7D7A787572706D6B686563605E5B585653514E4B494644413E3C393734312F2C";
constant INIT_H_IANA_61 : bit_vector(255 downto 0) := X"1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F";
constant INIT_L_IANA_61 : bit_vector(255 downto 0) := X"D0CDCBC8C5C3C0BEBBB8B6B3B1AEABA9A6A4A19E9C999794918F8C8A8784827F";
constant INIT_H_IANA_62 : bit_vector(255 downto 0) := X"20202020202020202020202020201F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F";
constant INIT_L_IANA_62 : bit_vector(255 downto 0) := X"23201E1B191613110E0C09060401FFFCF9F7F4F2EFECEAE7E5E2DFDDDAD8D5D2";
constant INIT_H_IANA_63 : bit_vector(255 downto 0) := X"2020202020202020202020202020202020202020202020202020202020202020";
constant INIT_L_IANA_63 : bit_vector(255 downto 0) := X"7674716E6C696764615F5C5A5754524F4D4A474542403D3A383533302D2B2826";
constant INIT_H_IANA_64 : bit_vector(255 downto 0) := X"2020202020202020202020202020202020202020202020202020202020202020";
constant INIT_L_IANA_64 : bit_vector(255 downto 0) := X"C9C7C4C1BFBCBAB7B4B2AFADAAA7A5A2A09D9A989593908D8B888683807E7B79";
constant INIT_H_IANA_65 : bit_vector(255 downto 0) := X"2121212121212121212121212020202020202020202020202020202020202020";
constant INIT_L_IANA_65 : bit_vector(255 downto 0) := X"1C1A1715120F0D0A08050200FDFBF8F5F3F0EEEBE8E6E3E1DEDBD9D6D4D1CECC";
constant INIT_H_IANA_66 : bit_vector(255 downto 0) := X"2121212121212121212121212121212121212121212121212121212121212121";
constant INIT_L_IANA_66 : bit_vector(255 downto 0) := X"6F6D6A686563605D5B585653504E4B494643413E3C393634312F2C292724221F";
constant INIT_H_IANA_67 : bit_vector(255 downto 0) := X"2121212121212121212121212121212121212121212121212121212121212121";
constant INIT_L_IANA_67 : bit_vector(255 downto 0) := X"C3C0BDBBB8B6B3B0AEABA9A6A3A19E9C999694918F8C898784827F7C7A777572";
constant INIT_H_IANA_68 : bit_vector(255 downto 0) := X"2222222222222222222121212121212121212121212121212121212121212121";
constant INIT_L_IANA_68 : bit_vector(255 downto 0) := X"1613110E0B09060401FEFCF9F7F4F1EFECEAE7E4E2DFDDDAD7D5D2D0CDCAC8C5";
constant INIT_H_IANA_69 : bit_vector(255 downto 0) := X"2222222222222222222222222222222222222222222222222222222222222222";
constant INIT_L_IANA_69 : bit_vector(255 downto 0) := X"696664615F5C595754524F4C4A4745423F3D3A383532302D2B282523201E1B18";
constant INIT_H_IANA_6A : bit_vector(255 downto 0) := X"2222222222222222222222222222222222222222222222222222222222222222";
constant INIT_L_IANA_6A : bit_vector(255 downto 0) := X"BCB9B7B4B2AFACAAA7A5A29F9D9A989592908D8B888583807E7B787673716E6B";
constant INIT_H_IANA_6B : bit_vector(255 downto 0) := X"2323232323232322222222222222222222222222222222222222222222222222";
constant INIT_L_IANA_6B : bit_vector(255 downto 0) := X"0F0D0A07050200FDFAF8F5F3F0EDEBE8E6E3E0DEDBD9D6D3D1CECCC9C6C4C1BF";
constant INIT_H_IANA_6C : bit_vector(255 downto 0) := X"2323232323232323232323232323232323232323232323232323232323232323";
constant INIT_L_IANA_6C : bit_vector(255 downto 0) := X"62605D5A585553504E4B484643413E3B393634312E2C292724211F1C1A171412";
constant INIT_H_IANA_6D : bit_vector(255 downto 0) := X"2323232323232323232323232323232323232323232323232323232323232323";
constant INIT_L_IANA_6D : bit_vector(255 downto 0) := X"B5B3B0AEABA8A6A3A19E9B999694918E8C898784817F7C7A7774726F6D6A6765";
constant INIT_H_IANA_6E : bit_vector(255 downto 0) := X"2424242423232323232323232323232323232323232323232323232323232323";
constant INIT_L_IANA_6E : bit_vector(255 downto 0) := X"09060301FEFCF9F6F4F1EFECE9E7E4E2DFDCDAD7D5D2CFCDCAC8C5C2C0BDBBB8";
constant INIT_H_IANA_6F : bit_vector(255 downto 0) := X"2424242424242424242424242424242424242424242424242424242424242424";
constant INIT_L_IANA_6F : bit_vector(255 downto 0) := X"5C595654514F4C4A4744423F3D3A373532302D2A282523201D1B181613100E0B";
constant INIT_H_IANA_70 : bit_vector(255 downto 0) := X"2424242424242424242424242424242424242424242424242424242424242424";
constant INIT_L_IANA_70 : bit_vector(255 downto 0) := X"AFACAAA7A4A29F9D9A979592908D8A888583807D7B787673706E6B696663615E";
constant INIT_H_IANA_71 : bit_vector(255 downto 0) := X"2524242424242424242424242424242424242424242424242424242424242424";
constant INIT_L_IANA_71 : bit_vector(255 downto 0) := X"02FFFDFAF8F5F2F0EDEBE8E5E3E0DEDBD8D6D3D1CECBC9C6C4C1BEBCB9B7B4B1";
constant INIT_H_IANA_72 : bit_vector(255 downto 0) := X"2525252525252525252525252525252525252525252525252525252525252525";
constant INIT_L_IANA_72 : bit_vector(255 downto 0) := X"5552504D4B484543403E3B393633312E2C292624211F1C191714120F0C0A0705";
constant INIT_H_IANA_73 : bit_vector(255 downto 0) := X"2525252525252525252525252525252525252525252525252525252525252525";
constant INIT_L_IANA_73 : bit_vector(255 downto 0) := X"A8A6A3A09E9B999693918E8C898684817F7C797774726F6C6A6765625F5D5A58";
constant INIT_H_IANA_74 : bit_vector(255 downto 0) := X"2525252525252525252525252525252525252525252525252525252525252525";
constant INIT_L_IANA_74 : bit_vector(255 downto 0) := X"FBF9F6F4F1EEECE9E7E4E1DFDCDAD7D4D2CFCDCAC7C5C2C0BDBAB8B5B3B0ADAB";
constant INIT_H_IANA_75 : bit_vector(255 downto 0) := X"2626262626262626262626262626262626262626262626262626262626262625";
constant INIT_L_IANA_75 : bit_vector(255 downto 0) := X"4E4C494744413F3C3A3734322F2D2A282522201D1B181513100E0B08060301FE";
constant INIT_H_IANA_76 : bit_vector(255 downto 0) := X"2626262626262626262626262626262626262626262626262626262626262626";
constant INIT_L_IANA_76 : bit_vector(255 downto 0) := X"A29F9C9A9795928F8D8A888582807D7B787573706E6B686663615E5B59565451";
constant INIT_H_IANA_77 : bit_vector(255 downto 0) := X"2626262626262626262626262626262626262626262626262626262626262626";
constant INIT_L_IANA_77 : bit_vector(255 downto 0) := X"F5F2F0EDEAE8E5E3E0DDDBD8D6D3D0CECBC9C6C3C1BEBCB9B6B4B1AFACA9A7A4";
constant INIT_H_IANA_78 : bit_vector(255 downto 0) := X"2727272727272727272727272727272727272727272727272727272726262626";
constant INIT_L_IANA_78 : bit_vector(255 downto 0) := X"484543403D3B383633302E2B292624211E1C191714110F0C0A070402FFFDFAF7";
constant INIT_H_IANA_79 : bit_vector(255 downto 0) := X"2727272727272727272727272727272727272727272727272727272727272727";
constant INIT_L_IANA_79 : bit_vector(255 downto 0) := X"9B989693918E8B898684817E7C797774716F6C6A6764625F5D5A575552504D4A";
constant INIT_H_IANA_7A : bit_vector(255 downto 0) := X"2727272727272727272727272727272727272727272727272727272727272727";
constant INIT_L_IANA_7A : bit_vector(255 downto 0) := X"EEECE9E6E4E1DFDCD9D7D4D2CFCCCAC7C5C2BFBDBAB8B5B2B0ADABA8A5A3A09E";
constant INIT_H_IANA_7B : bit_vector(255 downto 0) := X"2828282828282828282828282828282828282828282828282828272727272727";
constant INIT_L_IANA_7B : bit_vector(255 downto 0) := X"413F3C393734322F2C2A2725221F1D1A181513100D0B08060300FEFBF9F6F3F1";
constant INIT_H_IANA_7C : bit_vector(255 downto 0) := X"2828282828282828282828282828282828282828282828282828282828282828";
constant INIT_L_IANA_7C : bit_vector(255 downto 0) := X"94928F8D8A878582807D7A787573706D6B686663605E5B595653514E4C494644";
constant INIT_H_IANA_7D : bit_vector(255 downto 0) := X"2828282828282828282828282828282828282828282828282828282828282828";
constant INIT_L_IANA_7D : bit_vector(255 downto 0) := X"E8E5E2E0DDDBD8D5D3D0CECBC8C6C3C1BEBBB9B6B4B1AEACA9A7A4A19F9C9A97";
constant INIT_H_IANA_7E : bit_vector(255 downto 0) := X"2929292929292929292929292929292929292929292929282828282828282828";
constant INIT_L_IANA_7E : bit_vector(255 downto 0) := X"3B383533302E2B282623211E1B191614110F0C09070402FFFCFAF7F5F2EFEDEA";
constant INIT_H_IANA_7F : bit_vector(255 downto 0) := X"2929292929292929292929292929292929292929292929292929292929292929";
constant INIT_L_IANA_7F : bit_vector(255 downto 0) := X"8E8B898683817E7C797674716F6C696764625F5C5A5755524F4D4A484542403D";
constant INIT_H_IDIG_00 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IDIG_00 : bit_vector(255 downto 0) := X"282625242321201F1D1C1B19181716141312100F0E0C0B0A0907060503020100";
constant INIT_H_IDIG_01 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IDIG_01 : bit_vector(255 downto 0) := X"51504F4D4C4B4A484746444342403F3E3D3B3A39373635333231302E2D2C2A29";
constant INIT_H_IDIG_02 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IDIG_02 : bit_vector(255 downto 0) := X"7B7A787776747372716F6E6D6B6A69676665646261605E5D5C5A595857555453";
constant INIT_H_IDIG_03 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IDIG_03 : bit_vector(255 downto 0) := X"A4A3A2A19F9E9D9B9A99979695949291908E8D8C8A89888785848381807F7D7C";
constant INIT_H_IDIG_04 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IDIG_04 : bit_vector(255 downto 0) := X"CECDCBCAC9C8C6C5C4C2C1C0BEBDBCBBB9B8B7B5B4B3B1B0AFAEACABAAA8A7A6";
constant INIT_H_IDIG_05 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IDIG_05 : bit_vector(255 downto 0) := X"F8F6F5F4F2F1F0EFEDECEBE9E8E7E5E4E3E2E0DFDEDCDBDAD8D7D6D5D3D2D1CF";
constant INIT_H_IDIG_06 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101000000000000";
constant INIT_L_IDIG_06 : bit_vector(255 downto 0) := X"21201F1D1C1B19181715141312100F0E0C0B0A08070605030201FFFEFDFBFAF9";
constant INIT_H_IDIG_07 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IDIG_07 : bit_vector(255 downto 0) := X"4B49484746444342403F3E3C3B3A393736353332312F2E2D2C2A292826252422";
constant INIT_H_IDIG_08 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IDIG_08 : bit_vector(255 downto 0) := X"747372706F6E6D6B6A69676665636261605E5D5C5A59585655545351504F4D4C";
constant INIT_H_IDIG_09 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IDIG_09 : bit_vector(255 downto 0) := X"9E9D9B9A99979695939291908E8D8C8A89888685848381807F7D7C7B79787776";
constant INIT_H_IDIG_0A : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IDIG_0A : bit_vector(255 downto 0) := X"C7C6C5C4C2C1C0BEBDBCBAB9B8B7B5B4B3B1B0AFADACABAAA8A7A6A4A3A2A09F";
constant INIT_H_IDIG_0B : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IDIG_0B : bit_vector(255 downto 0) := X"F1F0EEEDECEAE9E8E7E5E4E3E1E0DFDEDCDBDAD8D7D6D4D3D2D1CFCECDCBCAC9";
constant INIT_H_IDIG_0C : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020101010101010101010101";
constant INIT_L_IDIG_0C : bit_vector(255 downto 0) := X"1B19181715141311100F0E0C0B0A08070604030201FFFEFDFBFAF9F7F6F5F4F2";
constant INIT_H_IDIG_0D : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IDIG_0D : bit_vector(255 downto 0) := X"444342403F3E3C3B3A383736353332312F2E2D2B2A29282625242221201E1D1C";
constant INIT_H_IDIG_0E : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IDIG_0E : bit_vector(255 downto 0) := X"6E6C6B6A686766656362615F5E5D5C5A59585655545251504F4D4C4B49484745";
constant INIT_H_IDIG_0F : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IDIG_0F : bit_vector(255 downto 0) := X"9796959392918F8E8D8C8A89888685848281807F7D7C7B79787775747372706F";
constant INIT_H_IDIG_10 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IDIG_10 : bit_vector(255 downto 0) := X"C1C0BEBDBCBAB9B8B6B5B4B3B1B0AFADACABA9A8A7A6A4A3A2A09F9E9C9B9A99";
constant INIT_H_IDIG_11 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IDIG_11 : bit_vector(255 downto 0) := X"EAE9E8E6E5E4E3E1E0DFDDDCDBDAD8D7D6D4D3D2D0CFCECDCBCAC9C7C6C5C3C2";
constant INIT_H_IDIG_12 : bit_vector(255 downto 0) := X"0303030303030303030303030303030302020202020202020202020202020202";
constant INIT_L_IDIG_12 : bit_vector(255 downto 0) := X"141311100F0D0C0B0A08070604030200FFFEFDFBFAF9F7F6F5F3F2F1F0EEEDEC";
constant INIT_H_IDIG_13 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IDIG_13 : bit_vector(255 downto 0) := X"3E3C3B3A383736343332312F2E2D2B2A29272625242221201E1D1C1A19181715";
constant INIT_H_IDIG_14 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IDIG_14 : bit_vector(255 downto 0) := X"6766646362615F5E5D5B5A59575655545251504E4D4C4B49484745444341403F";
constant INIT_H_IDIG_15 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IDIG_15 : bit_vector(255 downto 0) := X"918F8E8D8B8A89888685848281807E7D7C7B79787775747371706F6E6C6B6A68";
constant INIT_H_IDIG_16 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IDIG_16 : bit_vector(255 downto 0) := X"BAB9B8B6B5B4B2B1B0AFADACABA9A8A7A5A4A3A2A09F9E9C9B9A989796959392";
constant INIT_H_IDIG_17 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IDIG_17 : bit_vector(255 downto 0) := X"E4E2E1E0DFDDDCDBD9D8D7D5D4D3D2D0CFCECCCBCAC9C7C6C5C3C2C1BFBEBDBC";
constant INIT_H_IDIG_18 : bit_vector(255 downto 0) := X"0404040404040404040404030303030303030303030303030303030303030303";
constant INIT_L_IDIG_18 : bit_vector(255 downto 0) := X"0D0C0B0908070604030200FFFEFCFBFAF9F7F6F5F3F2F1EFEEEDECEAE9E8E6E5";
constant INIT_H_IDIG_19 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IDIG_19 : bit_vector(255 downto 0) := X"3736343332302F2E2D2B2A29272625232221201E1D1C1A19181615141311100F";
constant INIT_H_IDIG_1A : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IDIG_1A : bit_vector(255 downto 0) := X"605F5E5D5B5A59575655535251504E4D4C4A49484745444341403F3D3C3B3A38";
constant INIT_H_IDIG_1B : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IDIG_1B : bit_vector(255 downto 0) := X"8A89878685848281807E7D7C7A79787775747371706F6D6C6B6A686766646362";
constant INIT_H_IDIG_1C : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IDIG_1C : bit_vector(255 downto 0) := X"B4B2B1B0AEADACABA9A8A7A5A4A3A1A09F9E9C9B9A989796949392918F8E8D8B";
constant INIT_H_IDIG_1D : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IDIG_1D : bit_vector(255 downto 0) := X"DDDCDBD9D8D7D5D4D3D1D0CFCECCCBCAC8C7C6C5C3C2C1BFBEBDBBBAB9B8B6B5";
constant INIT_H_IDIG_1E : bit_vector(255 downto 0) := X"0505050505050404040404040404040404040404040404040404040404040404";
constant INIT_L_IDIG_1E : bit_vector(255 downto 0) := X"070504030200FFFEFCFBFAF8F7F6F5F3F2F1EFEEEDEBEAE9E8E6E5E4E2E1E0DE";
constant INIT_H_IDIG_1F : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IDIG_1F : bit_vector(255 downto 0) := X"302F2E2C2B2A292726252322211F1E1D1C1A19181615141211100F0D0C0B0908";
constant INIT_H_IDIG_20 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IDIG_20 : bit_vector(255 downto 0) := X"5A595756555352514F4E4D4C4A49484645444241403F3D3C3B39383736343332";
constant INIT_H_IDIG_21 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IDIG_21 : bit_vector(255 downto 0) := X"838281807E7D7C7A79787675747371706F6D6C6B69686766646362605F5E5C5B";
constant INIT_H_IDIG_22 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IDIG_22 : bit_vector(255 downto 0) := X"ADACAAA9A8A7A5A4A3A1A09F9D9C9B9A989796949392908F8E8D8B8A89878685";
constant INIT_H_IDIG_23 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IDIG_23 : bit_vector(255 downto 0) := X"D7D5D4D3D1D0CFCDCCCBCAC8C7C6C4C3C2C0BFBEBDBBBAB9B7B6B5B4B2B1B0AE";
constant INIT_H_IDIG_24 : bit_vector(255 downto 0) := X"0605050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IDIG_24 : bit_vector(255 downto 0) := X"00FFFEFCFBFAF8F7F6F4F3F2F1EFEEEDEBEAE9E7E6E5E4E2E1E0DEDDDCDAD9D8";
constant INIT_H_IDIG_25 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IDIG_25 : bit_vector(255 downto 0) := X"2A282726252322211F1E1D1B1A19181615141211100E0D0C0B09080705040301";
constant INIT_H_IDIG_26 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IDIG_26 : bit_vector(255 downto 0) := X"5352514F4E4D4B4A49484645444241403E3D3C3B39383735343332302F2E2C2B";
constant INIT_H_IDIG_27 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IDIG_27 : bit_vector(255 downto 0) := X"7D7C7A79787675747271706F6D6C6B69686765646362605F5E5C5B5A58575655";
constant INIT_H_IDIG_28 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IDIG_28 : bit_vector(255 downto 0) := X"A6A5A4A3A1A09F9D9C9B99989796949392908F8E8C8B8A898786858382817F7E";
constant INIT_H_IDIG_29 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IDIG_29 : bit_vector(255 downto 0) := X"D0CFCDCCCBC9C8C7C6C4C3C2C0BFBEBCBBBAB9B7B6B5B3B2B1AFAEADACAAA9A8";
constant INIT_H_IDIG_2A : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IDIG_2A : bit_vector(255 downto 0) := X"FAF8F7F6F4F3F2F0EFEEEDEBEAE9E7E6E5E3E2E1E0DEDDDCDAD9D8D6D5D4D3D1";
constant INIT_H_IDIG_2B : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070706060606";
constant INIT_L_IDIG_2B : bit_vector(255 downto 0) := X"2322211F1E1D1B1A19171615141211100E0D0C0A0908070504030100FFFDFCFB";
constant INIT_H_IDIG_2C : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IDIG_2C : bit_vector(255 downto 0) := X"4D4B4A49474645444241403E3D3C3A39383735343331302F2D2C2B2A28272624";
constant INIT_H_IDIG_2D : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IDIG_2D : bit_vector(255 downto 0) := X"7675747271706E6D6C6B69686765646361605F5E5C5B5A585756545352514F4E";
constant INIT_H_IDIG_2E : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IDIG_2E : bit_vector(255 downto 0) := X"A09F9D9C9B99989795949392908F8E8C8B8A888786858382817F7E7D7B7A7978";
constant INIT_H_IDIG_2F : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IDIG_2F : bit_vector(255 downto 0) := X"C9C8C7C5C4C3C2C0BFBEBCBBBAB8B7B6B5B3B2B1AFAEADABAAA9A8A6A5A4A2A1";
constant INIT_H_IDIG_30 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IDIG_30 : bit_vector(255 downto 0) := X"F3F2F0EFEEECEBEAE9E7E6E5E3E2E1DFDEDDDCDAD9D8D6D5D4D2D1D0CFCDCCCB";
constant INIT_H_IDIG_31 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808070707070707070707";
constant INIT_L_IDIG_31 : bit_vector(255 downto 0) := X"1D1B1A19171615131211100E0D0C0A0908060504030100FFFDFCFBF9F8F7F6F4";
constant INIT_H_IDIG_32 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IDIG_32 : bit_vector(255 downto 0) := X"4645434241403E3D3C3A39383635343331302F2D2C2B29282726242322201F1E";
constant INIT_H_IDIG_33 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IDIG_33 : bit_vector(255 downto 0) := X"706E6D6C6A69686765646361605F5D5C5B5A585756545352504F4E4D4B4A4947";
constant INIT_H_IDIG_34 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IDIG_34 : bit_vector(255 downto 0) := X"99989795949391908F8E8C8B8A888786848382817F7E7D7B7A79777675747271";
constant INIT_H_IDIG_35 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IDIG_35 : bit_vector(255 downto 0) := X"C3C1C0BFBEBCBBBAB8B7B6B4B3B2B1AFAEADABAAA9A7A6A5A4A2A1A09E9D9C9A";
constant INIT_H_IDIG_36 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IDIG_36 : bit_vector(255 downto 0) := X"ECEBEAE8E7E6E5E3E2E1DFDEDDDBDAD9D8D6D5D4D2D1D0CECDCCCBC9C8C7C5C4";
constant INIT_H_IDIG_37 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090808080808080808080808080808";
constant INIT_L_IDIG_37 : bit_vector(255 downto 0) := X"16151312110F0E0D0C0A0908060504020100FFFDFCFBF9F8F7F5F4F3F2F0EFEE";
constant INIT_H_IDIG_38 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IDIG_38 : bit_vector(255 downto 0) := X"3F3E3D3C3A39383635343231302F2D2C2B29282725242322201F1E1C1B1A1817";
constant INIT_H_IDIG_39 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IDIG_39 : bit_vector(255 downto 0) := X"69686665646361605F5D5C5B59585756545352504F4E4C4B4A49474645434241";
constant INIT_H_IDIG_3A : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IDIG_3A : bit_vector(255 downto 0) := X"9391908F8D8C8B8A888786848382807F7E7D7B7A79777675737271706E6D6C6A";
constant INIT_H_IDIG_3B : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IDIG_3B : bit_vector(255 downto 0) := X"BCBBBAB8B7B6B4B3B2B0AFAEADABAAA9A7A6A5A3A2A1A09E9D9C9A9998969594";
constant INIT_H_IDIG_3C : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IDIG_3C : bit_vector(255 downto 0) := X"E6E4E3E2E1DFDEDDDBDAD9D7D6D5D4D2D1D0CECDCCCAC9C8C7C5C4C3C1C0BFBD";
constant INIT_H_IDIG_3D : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A09090909090909090909090909090909090909";
constant INIT_L_IDIG_3D : bit_vector(255 downto 0) := X"0F0E0D0B0A0907060504020100FEFDFCFBF9F8F7F5F4F3F1F0EFEEECEBEAE8E7";
constant INIT_H_IDIG_3E : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_IDIG_3E : bit_vector(255 downto 0) := X"39383635343231302E2D2C2B29282725242321201F1E1C1B1A18171614131211";
constant INIT_H_IDIG_3F : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_IDIG_3F : bit_vector(255 downto 0) := X"6261605F5D5C5B59585755545352504F4E4C4B4A484746454342413F3E3D3B3A";
constant INIT_H_IDIG_40 : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_IDIG_40 : bit_vector(255 downto 0) := X"8C8B89888785848382807F7E7C7B7A797776757372716F6E6D6C6A6968666564";
constant INIT_H_IDIG_41 : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_IDIG_41 : bit_vector(255 downto 0) := X"B6B4B3B2B0AFAEACABAAA9A7A6A5A3A2A19F9E9D9C9A99989695949291908F8D";
constant INIT_H_IDIG_42 : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_IDIG_42 : bit_vector(255 downto 0) := X"DFDEDDDBDAD9D7D6D5D3D2D1D0CECDCCCAC9C8C6C5C4C3C1C0BFBDBCBBB9B8B7";
constant INIT_H_IDIG_43 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_IDIG_43 : bit_vector(255 downto 0) := X"0907060503020100FEFDFCFAF9F8F7F5F4F3F1F0EFEDECEBEAE8E7E6E4E3E2E0";
constant INIT_H_IDIG_44 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_IDIG_44 : bit_vector(255 downto 0) := X"3231302E2D2C2A29282725242321201F1D1C1B1A181716141312100F0E0D0B0A";
constant INIT_H_IDIG_45 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_IDIG_45 : bit_vector(255 downto 0) := X"5C5B59585755545351504F4E4C4B4A484746444342413F3E3D3B3A3937363534";
constant INIT_H_IDIG_46 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_IDIG_46 : bit_vector(255 downto 0) := X"85848381807F7E7C7B7A787776747372716F6E6D6B6A69686665646261605E5D";
constant INIT_H_IDIG_47 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_IDIG_47 : bit_vector(255 downto 0) := X"AFAEACABAAA8A7A6A5A3A2A19F9E9D9B9A99989695949291908E8D8C8B898887";
constant INIT_H_IDIG_48 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_IDIG_48 : bit_vector(255 downto 0) := X"D9D7D6D5D3D2D1CFCECDCCCAC9C8C6C5C4C2C1C0BFBDBCBBB9B8B7B5B4B3B2B0";
constant INIT_H_IDIG_49 : bit_vector(255 downto 0) := X"0C0C0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_IDIG_49 : bit_vector(255 downto 0) := X"0201FFFEFDFCFAF9F8F6F5F4F2F1F0EFEDECEBE9E8E7E6E4E3E2E0DFDEDCDBDA";
constant INIT_H_IDIG_4A : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_IDIG_4A : bit_vector(255 downto 0) := X"2C2A29282625242321201F1D1C1B19181716141312100F0E0C0B0A0907060503";
constant INIT_H_IDIG_4B : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_IDIG_4B : bit_vector(255 downto 0) := X"55545351504F4D4C4B4A484746444342403F3E3D3B3A39373635333231302E2D";
constant INIT_H_IDIG_4C : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_IDIG_4C : bit_vector(255 downto 0) := X"7F7D7C7B7A787776747372706F6E6D6B6A69676665646261605E5D5C5A595857";
constant INIT_H_IDIG_4D : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_IDIG_4D : bit_vector(255 downto 0) := X"A8A7A6A4A3A2A19F9E9D9B9A99979695949291908E8D8C8A8988878584838180";
constant INIT_H_IDIG_4E : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_IDIG_4E : bit_vector(255 downto 0) := X"D2D1CFCECDCBCAC9C8C6C5C4C2C1C0BEBDBCBBB9B8B7B5B4B3B1B0AFAEACABAA";
constant INIT_H_IDIG_4F : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_IDIG_4F : bit_vector(255 downto 0) := X"FBFAF9F8F6F5F4F2F1F0EEEDECEBE9E8E7E5E4E3E2E0DFDEDCDBDAD8D7D6D5D3";
constant INIT_H_IDIG_50 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0C0C0C";
constant INIT_L_IDIG_50 : bit_vector(255 downto 0) := X"25242221201F1D1C1B19181715141312100F0E0C0B0A08070605030201FFFEFD";
constant INIT_H_IDIG_51 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_IDIG_51 : bit_vector(255 downto 0) := X"4F4D4C4B49484746444342403F3E3C3B3A393736353332312F2E2D2C2A292826";
constant INIT_H_IDIG_52 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_IDIG_52 : bit_vector(255 downto 0) := X"787776747372706F6E6C6B6A696766656362615F5E5D5C5A5958565554535150";
constant INIT_H_IDIG_53 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_IDIG_53 : bit_vector(255 downto 0) := X"A2A09F9E9D9B9A99979695939291908E8D8C8A89888685848381807F7D7C7B79";
constant INIT_H_IDIG_54 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_IDIG_54 : bit_vector(255 downto 0) := X"CBCAC9C7C6C5C4C2C1C0BEBDBCBAB9B8B7B5B4B3B1B0AFADACABAAA8A7A6A4A3";
constant INIT_H_IDIG_55 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_IDIG_55 : bit_vector(255 downto 0) := X"F5F4F2F1F0EEEDECEAE9E8E7E5E4E3E1E0DFDDDCDBDAD8D7D6D4D3D2D1CFCECD";
constant INIT_H_IDIG_56 : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0D0D0D0D0D0D0D0D";
constant INIT_L_IDIG_56 : bit_vector(255 downto 0) := X"1E1D1C1B19181715141311100F0E0C0B0A08070604030201FFFEFDFBFAF9F7F6";
constant INIT_H_IDIG_57 : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_IDIG_57 : bit_vector(255 downto 0) := X"484745444342403F3E3C3B3A383736353332312F2E2D2B2A2928262524222120";
constant INIT_H_IDIG_58 : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_IDIG_58 : bit_vector(255 downto 0) := X"72706F6E6C6B6A686766656362615F5E5D5B5A59585655545251504F4D4C4B49";
constant INIT_H_IDIG_59 : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_IDIG_59 : bit_vector(255 downto 0) := X"9B9A999796959392918F8E8D8C8A89888685848281807F7D7C7B797877757473";
constant INIT_H_IDIG_5A : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_IDIG_5A : bit_vector(255 downto 0) := X"C5C3C2C1C0BEBDBCBAB9B8B6B5B4B3B1B0AFADACABA9A8A7A6A4A3A2A09F9E9C";
constant INIT_H_IDIG_5B : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_IDIG_5B : bit_vector(255 downto 0) := X"EEEDECEAE9E8E6E5E4E3E1E0DFDDDCDBD9D8D7D6D4D3D2D0CFCECCCBCAC9C7C6";
constant INIT_H_IDIG_5C : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_IDIG_5C : bit_vector(255 downto 0) := X"181715141311100F0D0C0B0A08070604030200FFFEFDFBFAF9F7F6F5F3F2F1F0";
constant INIT_H_IDIG_5D : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_IDIG_5D : bit_vector(255 downto 0) := X"41403F3E3C3B3A383736343332312F2E2D2B2A29272625242221201E1D1C1A19";
constant INIT_H_IDIG_5E : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_IDIG_5E : bit_vector(255 downto 0) := X"6B6A686766646362615F5E5D5B5A59575655545251504E4D4C4A494847454443";
constant INIT_H_IDIG_5F : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_IDIG_5F : bit_vector(255 downto 0) := X"959392918F8E8D8B8A89888685848281807E7D7C7B79787775747371706F6E6C";
constant INIT_H_IDIG_60 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_IDIG_60 : bit_vector(255 downto 0) := X"BEBDBCBAB9B8B6B5B4B2B1B0AFADACABA9A8A7A5A4A3A2A09F9E9C9B9A989796";
constant INIT_H_IDIG_61 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_IDIG_61 : bit_vector(255 downto 0) := X"E8E6E5E4E2E1E0DFDDDCDBD9D8D7D5D4D3D2D0CFCECCCBCAC8C7C6C5C3C2C1BF";
constant INIT_H_IDIG_62 : bit_vector(255 downto 0) := X"10101010101010101010101010100F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_IDIG_62 : bit_vector(255 downto 0) := X"11100F0D0C0B0908070604030200FFFEFCFBFAF9F7F6F5F3F2F1EFEEEDECEAE9";
constant INIT_H_IDIG_63 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_IDIG_63 : bit_vector(255 downto 0) := X"3B3A383736343332302F2E2D2B2A29272625232221201E1D1C1A191816151413";
constant INIT_H_IDIG_64 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_IDIG_64 : bit_vector(255 downto 0) := X"646362605F5E5D5B5A59575655535251504E4D4C4A49484645444341403F3D3C";
constant INIT_H_IDIG_65 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_IDIG_65 : bit_vector(255 downto 0) := X"8E8D8B8A89878685848281807E7D7C7A79787775747371706F6D6C6B6A686766";
constant INIT_H_IDIG_66 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_IDIG_66 : bit_vector(255 downto 0) := X"B7B6B5B4B2B1B0AEADACABA9A8A7A5A4A3A1A09F9E9C9B9A989796949392918F";
constant INIT_H_IDIG_67 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_IDIG_67 : bit_vector(255 downto 0) := X"E1E0DEDDDCDBD9D8D7D5D4D3D1D0CFCECCCBCAC8C7C6C4C3C2C1BFBEBDBBBAB9";
constant INIT_H_IDIG_68 : bit_vector(255 downto 0) := X"1111111111111111111010101010101010101010101010101010101010101010";
constant INIT_L_IDIG_68 : bit_vector(255 downto 0) := X"0B0908070504030200FFFEFCFBFAF8F7F6F5F3F2F1EFEEEDEBEAE9E8E6E5E4E2";
constant INIT_H_IDIG_69 : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_IDIG_69 : bit_vector(255 downto 0) := X"343332302F2E2C2B2A292726252322211F1E1D1C1A19181615141211100F0D0C";
constant INIT_H_IDIG_6A : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_IDIG_6A : bit_vector(255 downto 0) := X"5E5C5B5A595756555352514F4E4D4C4A49484645444241403F3D3C3B39383735";
constant INIT_H_IDIG_6B : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_IDIG_6B : bit_vector(255 downto 0) := X"878685838281807E7D7C7A79787675747371706F6D6C6B69686766646362605F";
constant INIT_H_IDIG_6C : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_IDIG_6C : bit_vector(255 downto 0) := X"B1B0AEADACAAA9A8A7A5A4A3A1A09F9D9C9B9A989796949392908F8E8D8B8A89";
constant INIT_H_IDIG_6D : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_IDIG_6D : bit_vector(255 downto 0) := X"DAD9D8D7D5D4D3D1D0CFCDCCCBCAC8C7C6C4C3C2C0BFBEBDBBBAB9B7B6B5B3B2";
constant INIT_H_IDIG_6E : bit_vector(255 downto 0) := X"1212121211111111111111111111111111111111111111111111111111111111";
constant INIT_L_IDIG_6E : bit_vector(255 downto 0) := X"04030100FFFEFCFBFAF8F7F6F4F3F2F1EFEEEDEBEAE9E7E6E5E4E2E1E0DEDDDC";
constant INIT_H_IDIG_6F : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_IDIG_6F : bit_vector(255 downto 0) := X"2E2C2B2A282726242322211F1E1D1B1A19181615141211100E0D0C0B09080705";
constant INIT_H_IDIG_70 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_IDIG_70 : bit_vector(255 downto 0) := X"5756555352514F4E4D4B4A49484645444241403E3D3C3B39383735343331302F";
constant INIT_H_IDIG_71 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_IDIG_71 : bit_vector(255 downto 0) := X"817F7E7D7C7A79787675747271706F6D6C6B69686765646362605F5E5C5B5A58";
constant INIT_H_IDIG_72 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_IDIG_72 : bit_vector(255 downto 0) := X"AAA9A8A6A5A4A2A1A09F9D9C9B99989796949392908F8E8C8B8A898786858382";
constant INIT_H_IDIG_73 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_IDIG_73 : bit_vector(255 downto 0) := X"D4D3D1D0CFCDCCCBC9C8C7C6C4C3C2C0BFBEBCBBBAB9B7B6B5B3B2B1AFAEADAC";
constant INIT_H_IDIG_74 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_IDIG_74 : bit_vector(255 downto 0) := X"FDFCFBFAF8F7F6F4F3F2F0EFEEEDEBEAE9E7E6E5E3E2E1E0DEDDDCDAD9D8D6D5";
constant INIT_H_IDIG_75 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131312";
constant INIT_L_IDIG_75 : bit_vector(255 downto 0) := X"2726242322201F1E1D1B1A19171615141211100E0D0C0A0908070504030100FF";
constant INIT_H_IDIG_76 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_IDIG_76 : bit_vector(255 downto 0) := X"514F4E4D4B4A49474645444241403E3D3C3A39383735343331302F2D2C2B2A28";
constant INIT_H_IDIG_77 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_IDIG_77 : bit_vector(255 downto 0) := X"7A79787675747271706E6D6C6B69686765646361605F5E5C5B5A585756545352";
constant INIT_H_IDIG_78 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_IDIG_78 : bit_vector(255 downto 0) := X"A4A2A1A09E9D9C9B99989795949392908F8E8C8B8A888786858382817F7E7D7B";
constant INIT_H_IDIG_79 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_IDIG_79 : bit_vector(255 downto 0) := X"CDCCCBC9C8C7C5C4C3C2C0BFBEBCBBBAB8B7B6B5B3B2B1AFAEADABAAA9A8A6A5";
constant INIT_H_IDIG_7A : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_IDIG_7A : bit_vector(255 downto 0) := X"F7F6F4F3F2F0EFEEECEBEAE9E7E6E5E3E2E1DFDEDDDCDAD9D8D6D5D4D2D1D0CF";
constant INIT_H_IDIG_7B : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414131313131313";
constant INIT_L_IDIG_7B : bit_vector(255 downto 0) := X"201F1E1C1B1A191716151312110F0E0D0C0A0908060504030100FFFDFCFBF9F8";
constant INIT_H_IDIG_7C : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_IDIG_7C : bit_vector(255 downto 0) := X"4A49474645434241403E3D3C3A39383635343331302F2D2C2B29282726242322";
constant INIT_H_IDIG_7D : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_IDIG_7D : bit_vector(255 downto 0) := X"747271706E6D6C6A69686765646361605F5D5C5B5A585756545352504F4E4D4B";
constant INIT_H_IDIG_7E : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_IDIG_7E : bit_vector(255 downto 0) := X"9D9C9A99989795949391908F8D8C8B8A888786848382817F7E7D7B7A79777675";
constant INIT_H_IDIG_7F : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_IDIG_7F : bit_vector(255 downto 0) := X"C7C5C4C3C1C0BFBEBCBBBAB8B7B6B4B3B2B1AFAEADABAAA9A7A6A5A4A2A1A09E";
constant INIT_H_IGUA_00 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_00 : bit_vector(255 downto 0) := X"12121111100F0F0E0E0D0C0C0B0A0A0909080707060605040403030201010000";
constant INIT_H_IGUA_01 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_01 : bit_vector(255 downto 0) := X"26252524242322222120201F1F1E1D1D1C1C1B1A1A1919181717161515141413";
constant INIT_H_IGUA_02 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_02 : bit_vector(255 downto 0) := X"39393838373636353534333332323130302F2F2E2D2D2C2B2B2A2A2928282727";
constant INIT_H_IGUA_03 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_03 : bit_vector(255 downto 0) := X"4D4C4C4B4B4A49494848474646454444434342414140403F3E3E3D3D3C3B3B3A";
constant INIT_H_IGUA_04 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_04 : bit_vector(255 downto 0) := X"61605F5F5E5E5D5C5C5B5A5A595958575756565554545353525151504F4F4E4E";
constant INIT_H_IGUA_05 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_05 : bit_vector(255 downto 0) := X"74737372727170706F6F6E6D6D6C6C6B6A6A6969686767666565646463626261";
constant INIT_H_IGUA_06 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_06 : bit_vector(255 downto 0) := X"88878686858584838382828180807F7E7E7D7D7C7B7B7A7A7978787777767575";
constant INIT_H_IGUA_07 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_07 : bit_vector(255 downto 0) := X"9B9B9A99999898979696959494939392919190908F8E8E8D8D8C8B8B8A898988";
constant INIT_H_IGUA_08 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_08 : bit_vector(255 downto 0) := X"AFAEADADACACABAAAAA9A9A8A7A7A6A6A5A4A4A3A3A2A1A1A09F9F9E9E9D9C9C";
constant INIT_H_IGUA_09 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_09 : bit_vector(255 downto 0) := X"C2C2C1C0C0BFBFBEBDBDBCBCBBBABAB9B8B8B7B7B6B5B5B4B4B3B2B2B1B1B0AF";
constant INIT_H_IGUA_0A : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_0A : bit_vector(255 downto 0) := X"D6D5D5D4D3D3D2D2D1D0D0CFCECECDCDCCCBCBCACAC9C8C8C7C7C6C5C5C4C3C3";
constant INIT_H_IGUA_0B : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_0B : bit_vector(255 downto 0) := X"E9E9E8E7E7E6E6E5E4E4E3E3E2E1E1E0E0DFDEDEDDDDDCDBDBDAD9D9D8D8D7D6";
constant INIT_H_IGUA_0C : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IGUA_0C : bit_vector(255 downto 0) := X"FDFCFCFBFAFAF9F9F8F7F7F6F6F5F4F4F3F2F2F1F1F0EFEFEEEEEDECECEBEBEA";
constant INIT_H_IGUA_0D : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010100000000";
constant INIT_L_IGUA_0D : bit_vector(255 downto 0) := X"10100F0F0E0D0D0C0C0B0A0A09080807070605050404030202010100FFFFFEFD";
constant INIT_H_IGUA_0E : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IGUA_0E : bit_vector(255 downto 0) := X"24232322212120201F1E1E1D1D1C1B1B1A1A1918181716161515141313121211";
constant INIT_H_IGUA_0F : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IGUA_0F : bit_vector(255 downto 0) := X"37373636353434333332313130302F2E2E2D2C2C2B2B2A292928282726262525";
constant INIT_H_IGUA_10 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IGUA_10 : bit_vector(255 downto 0) := X"4B4A4A494948474746464544444342424141403F3F3E3E3D3C3C3B3B3A393938";
constant INIT_H_IGUA_11 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IGUA_11 : bit_vector(255 downto 0) := X"5F5E5D5D5C5B5B5A5A595858575756555554545352525150504F4F4E4D4D4C4C";
constant INIT_H_IGUA_12 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IGUA_12 : bit_vector(255 downto 0) := X"72717170706F6E6E6D6D6C6B6B6A6A696868676666656564636362626160605F";
constant INIT_H_IGUA_13 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IGUA_13 : bit_vector(255 downto 0) := X"86858484838382818180807F7E7E7D7C7C7B7B7A797978787776767575747373";
constant INIT_H_IGUA_14 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IGUA_14 : bit_vector(255 downto 0) := X"999998979796959594949392929191908F8F8E8E8D8C8C8B8A8A898988878786";
constant INIT_H_IGUA_15 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IGUA_15 : bit_vector(255 downto 0) := X"ADACABABAAAAA9A8A8A7A7A6A5A5A4A4A3A2A2A1A0A09F9F9E9D9D9C9C9B9A9A";
constant INIT_H_IGUA_16 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IGUA_16 : bit_vector(255 downto 0) := X"C0C0BFBEBEBDBDBCBBBBBABAB9B8B8B7B6B6B5B5B4B3B3B2B2B1B0B0AFAFAEAD";
constant INIT_H_IGUA_17 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IGUA_17 : bit_vector(255 downto 0) := X"D4D3D3D2D1D1D0CFCFCECECDCCCCCBCBCAC9C9C8C8C7C6C6C5C4C4C3C3C2C1C1";
constant INIT_H_IGUA_18 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IGUA_18 : bit_vector(255 downto 0) := X"E7E7E6E5E5E4E4E3E2E2E1E1E0DFDFDEDEDDDCDCDBDADAD9D9D8D7D7D6D6D5D4";
constant INIT_H_IGUA_19 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IGUA_19 : bit_vector(255 downto 0) := X"FBFAFAF9F8F8F7F7F6F5F5F4F3F3F2F2F1F0F0EFEFEEEDEDECECEBEAEAE9E9E8";
constant INIT_H_IGUA_1A : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020201010101010101";
constant INIT_L_IGUA_1A : bit_vector(255 downto 0) := X"0E0E0D0D0C0B0B0A0909080807060605050403030202010000FFFEFEFDFDFCFB";
constant INIT_H_IGUA_1B : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IGUA_1B : bit_vector(255 downto 0) := X"222121201F1F1E1E1D1C1C1B1B1A19191818171616151414131312111110100F";
constant INIT_H_IGUA_1C : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IGUA_1C : bit_vector(255 downto 0) := X"353534343332323131302F2F2E2D2D2C2C2B2A2A292928272726262524242323";
constant INIT_H_IGUA_1D : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IGUA_1D : bit_vector(255 downto 0) := X"494848474746454544434342424140403F3F3E3D3D3C3C3B3A3A393838373736";
constant INIT_H_IGUA_1E : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IGUA_1E : bit_vector(255 downto 0) := X"5D5C5B5B5A59595858575656555554535352525150504F4E4E4D4D4C4B4B4A4A";
constant INIT_H_IGUA_1F : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IGUA_1F : bit_vector(255 downto 0) := X"706F6F6E6E6D6C6C6B6B6A69696867676666656464636362616160605F5E5E5D";
constant INIT_H_IGUA_20 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IGUA_20 : bit_vector(255 downto 0) := X"848382828181807F7F7E7D7D7C7C7B7A7A797978777776767574747372727171";
constant INIT_H_IGUA_21 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IGUA_21 : bit_vector(255 downto 0) := X"979796959594939392929190908F8F8E8D8D8C8C8B8A8A898888878786858584";
constant INIT_H_IGUA_22 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IGUA_22 : bit_vector(255 downto 0) := X"ABAAA9A9A8A8A7A6A6A5A5A4A3A3A2A1A1A0A09F9E9E9D9D9C9B9B9A9A999898";
constant INIT_H_IGUA_23 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IGUA_23 : bit_vector(255 downto 0) := X"BEBEBDBCBCBBBBBAB9B9B8B7B7B6B6B5B4B4B3B3B2B1B1B0B0AFAEAEADACACAB";
constant INIT_H_IGUA_24 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IGUA_24 : bit_vector(255 downto 0) := X"D2D1D1D0CFCFCECDCDCCCCCBCACAC9C9C8C7C7C6C6C5C4C4C3C2C2C1C1C0BFBF";
constant INIT_H_IGUA_25 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IGUA_25 : bit_vector(255 downto 0) := X"E5E5E4E3E3E2E2E1E0E0DFDFDEDDDDDCDBDBDADAD9D8D8D7D7D6D5D5D4D4D3D2";
constant INIT_H_IGUA_26 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IGUA_26 : bit_vector(255 downto 0) := X"F9F8F8F7F6F6F5F5F4F3F3F2F1F1F0F0EFEEEEEDEDECEBEBEAEAE9E8E8E7E6E6";
constant INIT_H_IGUA_27 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030302020202020202020202";
constant INIT_L_IGUA_27 : bit_vector(255 downto 0) := X"0C0C0B0A0A0909080707060605040403030201010000FFFEFEFDFCFCFBFBFAF9";
constant INIT_H_IGUA_28 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IGUA_28 : bit_vector(255 downto 0) := X"201F1F1E1D1D1C1C1B1A1A191918171716151514141312121111100F0F0E0E0D";
constant INIT_H_IGUA_29 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IGUA_29 : bit_vector(255 downto 0) := X"333332323130302F2F2E2D2D2C2B2B2A2A292828272726252524242322222120";
constant INIT_H_IGUA_2A : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IGUA_2A : bit_vector(255 downto 0) := X"474646454444434342414140403F3E3E3D3D3C3B3B3A3A393838373636353534";
constant INIT_H_IGUA_2B : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IGUA_2B : bit_vector(255 downto 0) := X"5A5A595958575756565554545353525151504F4F4E4E4D4C4C4B4B4A49494848";
constant INIT_H_IGUA_2C : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IGUA_2C : bit_vector(255 downto 0) := X"6E6D6D6C6C6B6A6A696968676766656564646362626161605F5F5E5E5D5C5C5B";
constant INIT_H_IGUA_2D : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IGUA_2D : bit_vector(255 downto 0) := X"828180807F7E7E7D7D7C7B7B7A7A797878777776757574747372727170706F6F";
constant INIT_H_IGUA_2E : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IGUA_2E : bit_vector(255 downto 0) := X"959494939392919190908F8E8E8D8D8C8B8B8A89898888878686858584838382";
constant INIT_H_IGUA_2F : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IGUA_2F : bit_vector(255 downto 0) := X"A9A8A7A7A6A6A5A4A4A3A3A2A1A1A09F9F9E9E9D9C9C9B9B9A99999898979696";
constant INIT_H_IGUA_30 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IGUA_30 : bit_vector(255 downto 0) := X"BCBCBBBABAB9B8B8B7B7B6B5B5B4B4B3B2B2B1B1B0AFAFAEAEADACACABAAAAA9";
constant INIT_H_IGUA_31 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IGUA_31 : bit_vector(255 downto 0) := X"D0CFCECECDCDCCCBCBCACAC9C8C8C7C7C6C5C5C4C3C3C2C2C1C0C0BFBFBEBDBD";
constant INIT_H_IGUA_32 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IGUA_32 : bit_vector(255 downto 0) := X"E3E3E2E1E1E0E0DFDEDEDDDDDCDBDBDAD9D9D8D8D7D6D6D5D5D4D3D3D2D2D1D0";
constant INIT_H_IGUA_33 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IGUA_33 : bit_vector(255 downto 0) := X"F7F6F6F5F4F4F3F2F2F1F1F0EFEFEEEEEDECECEBEBEAE9E9E8E7E7E6E6E5E4E4";
constant INIT_H_IGUA_34 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040303030303030303030303030303";
constant INIT_L_IGUA_34 : bit_vector(255 downto 0) := X"0A0A09080807070605050404030202010100FFFFFEFDFDFCFCFBFAFAF9F9F8F7";
constant INIT_H_IGUA_35 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IGUA_35 : bit_vector(255 downto 0) := X"1E1D1D1C1B1B1A1A191818171716151514131312121110100F0F0E0D0D0C0C0B";
constant INIT_H_IGUA_36 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IGUA_36 : bit_vector(255 downto 0) := X"313130302F2E2E2D2C2C2B2B2A29292828272626252524232322212120201F1E";
constant INIT_H_IGUA_37 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IGUA_37 : bit_vector(255 downto 0) := X"4544444342424141403F3F3E3E3D3C3C3B3B3A39393837373636353434333332";
constant INIT_H_IGUA_38 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IGUA_38 : bit_vector(255 downto 0) := X"5858575756555554545352525151504F4F4E4D4D4C4C4B4A4A49494847474646";
constant INIT_H_IGUA_39 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IGUA_39 : bit_vector(255 downto 0) := X"6C6B6B6A6A696868676666656564636362626160605F5F5E5D5D5C5B5B5A5A59";
constant INIT_H_IGUA_3A : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IGUA_3A : bit_vector(255 downto 0) := X"807F7E7E7D7C7C7B7B7A79797878777676757574737372717170706F6E6E6D6D";
constant INIT_H_IGUA_3B : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IGUA_3B : bit_vector(255 downto 0) := X"9392929191908F8F8E8E8D8C8C8B8B8A89898887878686858484838382818180";
constant INIT_H_IGUA_3C : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IGUA_3C : bit_vector(255 downto 0) := X"A7A6A5A5A4A4A3A2A2A1A0A09F9F9E9D9D9C9C9B9A9A99999897979695959494";
constant INIT_H_IGUA_3D : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IGUA_3D : bit_vector(255 downto 0) := X"BABAB9B8B8B7B6B6B5B5B4B3B3B2B2B1B0B0AFAFAEADADACABABAAAAA9A8A8A7";
constant INIT_H_IGUA_3E : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IGUA_3E : bit_vector(255 downto 0) := X"CECDCCCCCBCBCAC9C9C8C8C7C6C6C5C5C4C3C3C2C1C1C0C0BFBEBEBDBDBCBBBB";
constant INIT_H_IGUA_3F : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IGUA_3F : bit_vector(255 downto 0) := X"E1E1E0DFDFDEDEDDDCDCDBDADAD9D9D8D7D7D6D6D5D4D4D3D3D2D1D1D0CFCFCE";
constant INIT_H_IGUA_40 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IGUA_40 : bit_vector(255 downto 0) := X"F5F4F4F3F2F2F1F0F0EFEFEEEDEDECECEBEAEAE9E9E8E7E7E6E5E5E4E4E3E2E2";
constant INIT_H_IGUA_41 : bit_vector(255 downto 0) := X"0505050505050505050505050505050404040404040404040404040404040404";
constant INIT_L_IGUA_41 : bit_vector(255 downto 0) := X"080807060605050403030202010000FFFEFEFDFDFCFBFBFAFAF9F8F8F7F7F6F5";
constant INIT_H_IGUA_42 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IGUA_42 : bit_vector(255 downto 0) := X"1C1B1B1A19191818171616151414131312111110100F0E0E0D0D0C0B0B0A0909";
constant INIT_H_IGUA_43 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IGUA_43 : bit_vector(255 downto 0) := X"2F2F2E2E2D2C2C2B2A2A292928272726262524242323222121201F1F1E1E1D1C";
constant INIT_H_IGUA_44 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IGUA_44 : bit_vector(255 downto 0) := X"4342424140403F3F3E3D3D3C3C3B3A3A39383837373635353434333232313130";
constant INIT_H_IGUA_45 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IGUA_45 : bit_vector(255 downto 0) := X"5656555554535352525150504F4E4E4D4D4C4B4B4A4A49484847474645454443";
constant INIT_H_IGUA_46 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IGUA_46 : bit_vector(255 downto 0) := X"6A69696868676666656464636362616160605F5E5E5D5D5C5B5B5A5959585857";
constant INIT_H_IGUA_47 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IGUA_47 : bit_vector(255 downto 0) := X"7D7D7C7C7B7A7A797978777776767574747372727171706F6F6E6E6D6C6C6B6B";
constant INIT_H_IGUA_48 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IGUA_48 : bit_vector(255 downto 0) := X"9190908F8F8E8D8D8C8C8B8A8A898888878786858584848382828181807F7F7E";
constant INIT_H_IGUA_49 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IGUA_49 : bit_vector(255 downto 0) := X"A5A4A3A3A2A2A1A0A09F9E9E9D9D9C9B9B9A9A99989897979695959493939292";
constant INIT_H_IGUA_4A : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IGUA_4A : bit_vector(255 downto 0) := X"B8B7B7B6B6B5B4B4B3B3B2B1B1B0B0AFAEAEADACACABABAAA9A9A8A8A7A6A6A5";
constant INIT_H_IGUA_4B : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IGUA_4B : bit_vector(255 downto 0) := X"CCCBCACAC9C9C8C7C7C6C6C5C4C4C3C2C2C1C1C0BFBFBEBEBDBCBCBBBBBAB9B9";
constant INIT_H_IGUA_4C : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IGUA_4C : bit_vector(255 downto 0) := X"DFDFDEDDDDDCDBDBDADAD9D8D8D7D7D6D5D5D4D4D3D2D2D1D1D0CFCFCECDCDCC";
constant INIT_H_IGUA_4D : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IGUA_4D : bit_vector(255 downto 0) := X"F3F2F1F1F0F0EFEEEEEDEDECEBEBEAEAE9E8E8E7E6E6E5E5E4E3E3E2E2E1E0E0";
constant INIT_H_IGUA_4E : bit_vector(255 downto 0) := X"0606060606060606060606060505050505050505050505050505050505050505";
constant INIT_L_IGUA_4E : bit_vector(255 downto 0) := X"060605040403030201010000FFFEFEFDFCFCFBFBFAF9F9F8F8F7F6F6F5F5F4F3";
constant INIT_H_IGUA_4F : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_4F : bit_vector(255 downto 0) := X"1A191918171716151514141312121111100F0F0E0E0D0C0C0B0B0A0909080707";
constant INIT_H_IGUA_50 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_50 : bit_vector(255 downto 0) := X"2D2D2C2B2B2A2A292828272726252524242322222120201F1F1E1D1D1C1C1B1A";
constant INIT_H_IGUA_51 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_51 : bit_vector(255 downto 0) := X"4140403F3E3E3D3D3C3B3B3A3A393838373636353534333332323130302F2F2E";
constant INIT_H_IGUA_52 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_52 : bit_vector(255 downto 0) := X"54545353525151504F4F4E4E4D4C4C4B4B4A4949484847464645454443434241";
constant INIT_H_IGUA_53 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_53 : bit_vector(255 downto 0) := X"68676766656564646362626161605F5F5E5E5D5C5C5B5A5A5959585757565655";
constant INIT_H_IGUA_54 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_54 : bit_vector(255 downto 0) := X"7B7B7A7A797878777776757574747372727170706F6F6E6D6D6C6C6B6A6A6969";
constant INIT_H_IGUA_55 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_55 : bit_vector(255 downto 0) := X"8F8E8E8D8D8C8B8B8A89898888878686858584838382828180807F7F7E7D7D7C";
constant INIT_H_IGUA_56 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_56 : bit_vector(255 downto 0) := X"A3A2A1A1A09F9F9E9E9D9C9C9B9B9A9999989897969695949493939291919090";
constant INIT_H_IGUA_57 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_57 : bit_vector(255 downto 0) := X"B6B5B5B4B4B3B2B2B1B1B0AFAFAEAEADACACABAAAAA9A9A8A7A7A6A6A5A4A4A3";
constant INIT_H_IGUA_58 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_58 : bit_vector(255 downto 0) := X"CAC9C8C8C7C7C6C5C5C4C3C3C2C2C1C0C0BFBFBEBDBDBCBCBBBABAB9B8B8B7B7";
constant INIT_H_IGUA_59 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_59 : bit_vector(255 downto 0) := X"DDDDDCDBDBDAD9D9D8D8D7D6D6D5D5D4D3D3D2D2D1D0D0CFCECECDCDCCCBCBCA";
constant INIT_H_IGUA_5A : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_5A : bit_vector(255 downto 0) := X"F1F0EFEFEEEEEDECECEBEBEAE9E9E8E8E7E6E6E5E4E4E3E3E2E1E1E0E0DFDEDE";
constant INIT_H_IGUA_5B : bit_vector(255 downto 0) := X"0707070707070707060606060606060606060606060606060606060606060606";
constant INIT_L_IGUA_5B : bit_vector(255 downto 0) := X"0404030202010100FFFFFEFDFDFCFCFBFAFAF9F9F8F7F7F6F6F5F4F4F3F2F2F1";
constant INIT_H_IGUA_5C : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_5C : bit_vector(255 downto 0) := X"18171716151514131312121110100F0F0E0D0D0C0C0B0A0A0908080707060505";
constant INIT_H_IGUA_5D : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_5D : bit_vector(255 downto 0) := X"2B2B2A29292828272626252524232322222120201F1E1E1D1D1C1B1B1A1A1918";
constant INIT_H_IGUA_5E : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_5E : bit_vector(255 downto 0) := X"3F3E3E3D3C3C3B3B3A39393837373636353434333332313130302F2E2E2D2C2C";
constant INIT_H_IGUA_5F : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_5F : bit_vector(255 downto 0) := X"52525151504F4F4E4D4D4C4C4B4A4A494948474746464544444342424141403F";
constant INIT_H_IGUA_60 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_60 : bit_vector(255 downto 0) := X"66656564636362626160605F5F5E5D5D5C5C5B5A5A5958585757565555545453";
constant INIT_H_IGUA_61 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_61 : bit_vector(255 downto 0) := X"79797878777676757574737372717170706F6E6E6D6D6C6B6B6A6A6968686766";
constant INIT_H_IGUA_62 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_62 : bit_vector(255 downto 0) := X"8D8C8C8B8B8A89898887878686858484838382818180807F7E7E7D7C7C7B7B7A";
constant INIT_H_IGUA_63 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_63 : bit_vector(255 downto 0) := X"A0A09F9F9E9D9D9C9C9B9A9A999998979796969594949392929191908F8F8E8E";
constant INIT_H_IGUA_64 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_64 : bit_vector(255 downto 0) := X"B4B3B3B2B2B1B0B0AFAFAEADADACABABAAAAA9A8A8A7A7A6A5A5A4A4A3A2A2A1";
constant INIT_H_IGUA_65 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_65 : bit_vector(255 downto 0) := X"C8C7C6C6C5C5C4C3C3C2C1C1C0C0BFBEBEBDBDBCBBBBBABAB9B8B8B7B6B6B5B5";
constant INIT_H_IGUA_66 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_66 : bit_vector(255 downto 0) := X"DBDADAD9D9D8D7D7D6D6D5D4D4D3D3D2D1D1D0CFCFCECECDCCCCCBCBCAC9C9C8";
constant INIT_H_IGUA_67 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_67 : bit_vector(255 downto 0) := X"EFEEEDEDECECEBEAEAE9E9E8E7E7E6E5E5E4E4E3E2E2E1E1E0DFDFDEDEDDDCDC";
constant INIT_H_IGUA_68 : bit_vector(255 downto 0) := X"0808080808070707070707070707070707070707070707070707070707070707";
constant INIT_L_IGUA_68 : bit_vector(255 downto 0) := X"0202010000FFFFFEFDFDFCFBFBFAFAF9F8F8F7F7F6F5F5F4F4F3F2F2F1F0F0EF";
constant INIT_H_IGUA_69 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_69 : bit_vector(255 downto 0) := X"16151414131312111110100F0E0E0D0D0C0B0B0A090908080706060505040303";
constant INIT_H_IGUA_6A : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_6A : bit_vector(255 downto 0) := X"292928272726262524242323222121201F1F1E1E1D1C1C1B1B1A191918181716";
constant INIT_H_IGUA_6B : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_6B : bit_vector(255 downto 0) := X"3D3C3C3B3A3A393938373736353534343332323131302F2F2E2E2D2C2C2B2A2A";
constant INIT_H_IGUA_6C : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_6C : bit_vector(255 downto 0) := X"50504F4E4E4D4D4C4B4B4A4A494848474746454544434342424140403F3F3E3D";
constant INIT_H_IGUA_6D : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_6D : bit_vector(255 downto 0) := X"64636362616160605F5E5E5D5D5C5B5B5A595958585756565555545353525251";
constant INIT_H_IGUA_6E : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_6E : bit_vector(255 downto 0) := X"777776767574747373727171706F6F6E6E6D6C6C6B6B6A696968686766666564";
constant INIT_H_IGUA_6F : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_6F : bit_vector(255 downto 0) := X"8B8A8A898888878786858584848382828181807F7F7E7D7D7C7C7B7A7A797978";
constant INIT_H_IGUA_70 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_70 : bit_vector(255 downto 0) := X"9E9E9D9D9C9B9B9A9A999898979796959594939392929190908F8F8E8D8D8C8C";
constant INIT_H_IGUA_71 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_71 : bit_vector(255 downto 0) := X"B2B1B1B0B0AFAEAEADACACABABAAA9A9A8A8A7A6A6A5A5A4A3A3A2A2A1A0A09F";
constant INIT_H_IGUA_72 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_72 : bit_vector(255 downto 0) := X"C6C5C4C4C3C2C2C1C1C0BFBFBEBEBDBCBCBBBBBAB9B9B8B7B7B6B6B5B4B4B3B3";
constant INIT_H_IGUA_73 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_73 : bit_vector(255 downto 0) := X"D9D8D8D7D7D6D5D5D4D4D3D2D2D1D1D0CFCFCECDCDCCCCCBCACAC9C9C8C7C7C6";
constant INIT_H_IGUA_74 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_74 : bit_vector(255 downto 0) := X"EDECEBEBEAEAE9E8E8E7E6E6E5E5E4E3E3E2E2E1E0E0DFDFDEDDDDDCDCDBDADA";
constant INIT_H_IGUA_75 : bit_vector(255 downto 0) := X"0909080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IGUA_75 : bit_vector(255 downto 0) := X"0000FFFEFEFDFCFCFBFBFAF9F9F8F8F7F6F6F5F5F4F3F3F2F1F1F0F0EFEEEEED";
constant INIT_H_IGUA_76 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IGUA_76 : bit_vector(255 downto 0) := X"141312121111100F0F0E0E0D0C0C0B0B0A090908070706060504040303020101";
constant INIT_H_IGUA_77 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IGUA_77 : bit_vector(255 downto 0) := X"272726252524242322222120201F1F1E1D1D1C1C1B1A1A191918171716161514";
constant INIT_H_IGUA_78 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IGUA_78 : bit_vector(255 downto 0) := X"3B3A3A393838373636353534333332323130302F2F2E2D2D2C2B2B2A2A292828";
constant INIT_H_IGUA_79 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IGUA_79 : bit_vector(255 downto 0) := X"4E4E4D4C4C4B4B4A49494848474646454544434342414140403F3E3E3D3D3C3B";
constant INIT_H_IGUA_7A : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IGUA_7A : bit_vector(255 downto 0) := X"626161605F5F5E5E5D5C5C5B5A5A59595857575656555454535352515150504F";
constant INIT_H_IGUA_7B : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IGUA_7B : bit_vector(255 downto 0) := X"757574747372727170706F6F6E6D6D6C6C6B6A6A696968676766656564646362";
constant INIT_H_IGUA_7C : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IGUA_7C : bit_vector(255 downto 0) := X"898888878686858584838382828180807F7F7E7D7D7C7B7B7A7A797878777776";
constant INIT_H_IGUA_7D : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IGUA_7D : bit_vector(255 downto 0) := X"9C9C9B9B9A99999898979696959494939392919190908F8E8E8D8D8C8B8B8A8A";
constant INIT_H_IGUA_7E : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IGUA_7E : bit_vector(255 downto 0) := X"B0AFAFAEAEADACACABAAAAA9A9A8A7A7A6A6A5A4A4A3A3A2A1A1A09F9F9E9E9D";
constant INIT_H_IGUA_7F : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IGUA_7F : bit_vector(255 downto 0) := X"C3C3C2C2C1C0C0BFBFBEBDBDBCBCBBBABAB9B9B8B7B7B6B5B5B4B4B3B2B2B1B1";
constant INIT_H_IBIA_00 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IBIA_00 : bit_vector(255 downto 0) := X"5E5B5855524F4C494643403D393633302D2A2724211E1B1815120F0C09060300";
constant INIT_H_IBIA_01 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_IBIA_01 : bit_vector(255 downto 0) := X"C0BDBAB7B4B1ADAAA7A4A19E9B9895928F8C898683807D7A7773706D6A676461";
constant INIT_H_IBIA_02 : bit_vector(255 downto 0) := X"0101010101010101010101010000000000000000000000000000000000000000";
constant INIT_L_IBIA_02 : bit_vector(255 downto 0) := X"211E1B1815120F0C09060300FDFAF7F4F1EEEBE7E4E1DEDBD8D5D2CFCCC9C6C3";
constant INIT_H_IBIA_03 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IBIA_03 : bit_vector(255 downto 0) := X"83807D7A7774716E6B6865625F5B5855524F4C494643403D3A3734312E2B2825";
constant INIT_H_IBIA_04 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_IBIA_04 : bit_vector(255 downto 0) := X"E5E2DFDCD9D6D3CFCCC9C6C3C0BDBAB7B4B1AEABA8A5A29F9C9995928F8C8986";
constant INIT_H_IBIA_05 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020101010101010101";
constant INIT_L_IBIA_05 : bit_vector(255 downto 0) := X"4743403D3A3734312E2B2825221F1C191613100D09060300FDFAF7F4F1EEEBE8";
constant INIT_H_IBIA_06 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_IBIA_06 : bit_vector(255 downto 0) := X"A8A5A29F9C999693908D8A8784817D7A7774716E6B6865625F5C595653504D4A";
constant INIT_H_IBIA_07 : bit_vector(255 downto 0) := X"0303030302020202020202020202020202020202020202020202020202020202";
constant INIT_L_IBIA_07 : bit_vector(255 downto 0) := X"0A070401FEFBF8F5F1EEEBE8E5E2DFDCD9D6D3D0CDCAC7C4C1BEBBB7B4B1AEAB";
constant INIT_H_IBIA_08 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IBIA_08 : bit_vector(255 downto 0) := X"6C6965625F5C595653504D4A4744413E3B3835322F2B2825221F1C191613100D";
constant INIT_H_IBIA_09 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_IBIA_09 : bit_vector(255 downto 0) := X"CDCAC7C4C1BEBBB8B5B2AFACA9A6A39F9C999693908D8A8784817E7B7875726F";
constant INIT_H_IBIA_0A : bit_vector(255 downto 0) := X"0404040404040404040404040404040403030303030303030303030303030303";
constant INIT_L_IBIA_0A : bit_vector(255 downto 0) := X"2F2C292623201D1A1713100D0A070401FEFBF8F5F2EFECE9E6E3E0DDD9D6D3D0";
constant INIT_H_IBIA_0B : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IBIA_0B : bit_vector(255 downto 0) := X"918E8B8784817E7B7875726F6C696663605D5A5754514D4A4744413E3B383532";
constant INIT_H_IBIA_0C : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_IBIA_0C : bit_vector(255 downto 0) := X"F2EFECE9E6E3E0DDDAD7D4D1CECBC8C5C1BEBBB8B5B2AFACA9A6A3A09D9A9794";
constant INIT_H_IBIA_0D : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050504040404";
constant INIT_L_IBIA_0D : bit_vector(255 downto 0) := X"54514E4B4845423F3C3835322F2C292623201D1A1714110E0B080502FEFBF8F5";
constant INIT_H_IBIA_0E : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_IBIA_0E : bit_vector(255 downto 0) := X"B6B3B0ACA9A6A3A09D9A9794918E8B8885827F7C7976726F6C696663605D5A57";
constant INIT_H_IBIA_0F : bit_vector(255 downto 0) := X"0606060606060606050505050505050505050505050505050505050505050505";
constant INIT_L_IBIA_0F : bit_vector(255 downto 0) := X"1714110E0B080502FFFCF9F6F3F0EDEAE6E3E0DDDAD7D4D1CECBC8C5C2BFBCB9";
constant INIT_H_IBIA_10 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IBIA_10 : bit_vector(255 downto 0) := X"797673706D6A6764615E5A5754514E4B4845423F3C393633302D2A2724201D1A";
constant INIT_H_IBIA_11 : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_IBIA_11 : bit_vector(255 downto 0) := X"DBD8D5D2CECBC8C5C2BFBCB9B6B3B0ADAAA7A4A19E9B9894918E8B8885827F7C";
constant INIT_H_IBIA_12 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707060606060606060606060606";
constant INIT_L_IBIA_12 : bit_vector(255 downto 0) := X"3C393633302D2A2724211E1B1815120F0C080502FFFCF9F6F3F0EDEAE7E4E1DE";
constant INIT_H_IBIA_13 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IBIA_13 : bit_vector(255 downto 0) := X"9E9B9895928F8C898683807C797673706D6A6764615E5B5855524F4C4946423F";
constant INIT_H_IBIA_14 : bit_vector(255 downto 0) := X"0807070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_IBIA_14 : bit_vector(255 downto 0) := X"00FDFAF7F4F0EDEAE7E4E1DEDBD8D5D2CFCCC9C6C3C0BDBAB6B3B0ADAAA7A4A1";
constant INIT_H_IBIA_15 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IBIA_15 : bit_vector(255 downto 0) := X"615E5B5855524F4C494643403D3A3734312E2A2724211E1B1815120F0C090603";
constant INIT_H_IBIA_16 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_IBIA_16 : bit_vector(255 downto 0) := X"C3C0BDBAB7B4B1AEABA8A5A29E9B9895928F8C898683807D7A7774716E6B6864";
constant INIT_H_IBIA_17 : bit_vector(255 downto 0) := X"0909090909090909090909090908080808080808080808080808080808080808";
constant INIT_L_IBIA_17 : bit_vector(255 downto 0) := X"25221F1C1916120F0C09060300FDFAF7F4F1EEEBE8E5E2DFDCD8D5D2CFCCC9C6";
constant INIT_H_IBIA_18 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IBIA_18 : bit_vector(255 downto 0) := X"8683807D7A7774716E6B6865625F5C595653504C494643403D3A3734312E2B28";
constant INIT_H_IBIA_19 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_IBIA_19 : bit_vector(255 downto 0) := X"E8E5E2DFDCD9D6D3D0CDCAC7C3C0BDBAB7B4B1AEABA8A5A29F9C999693908D8A";
constant INIT_H_IBIA_1A : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A09090909090909";
constant INIT_L_IBIA_1A : bit_vector(255 downto 0) := X"4A4744413E3B3734312E2B2825221F1C191613100D0A070401FDFAF7F4F1EEEB";
constant INIT_H_IBIA_1B : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_IBIA_1B : bit_vector(255 downto 0) := X"ABA8A5A29F9C999693908D8A8784817E7B7875716E6B6865625F5C595653504D";
constant INIT_H_IBIA_1C : bit_vector(255 downto 0) := X"0B0B0B0B0B0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_IBIA_1C : bit_vector(255 downto 0) := X"0D0A070401FEFBF8F5F2EFECE9E5E2DFDCD9D6D3D0CDCAC7C4C1BEBBB8B5B2AF";
constant INIT_H_IBIA_1D : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_IBIA_1D : bit_vector(255 downto 0) := X"6F6C696663605D595653504D4A4744413E3B3835322F2C2926231F1C19161310";
constant INIT_H_IBIA_1E : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_IBIA_1E : bit_vector(255 downto 0) := X"D1CDCAC7C4C1BEBBB8B5B2AFACA9A6A3A09D9A9793908D8A8784817E7B787572";
constant INIT_H_IBIA_1F : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_IBIA_1F : bit_vector(255 downto 0) := X"322F2C292623201D1A1714110E0B070401FEFBF8F5F2EFECE9E6E3E0DDDAD7D4";
constant INIT_H_IBIA_20 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_IBIA_20 : bit_vector(255 downto 0) := X"94918E8B8885827F7B7875726F6C696663605D5A5754514E4B4845413E3B3835";
constant INIT_H_IBIA_21 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_IBIA_21 : bit_vector(255 downto 0) := X"F6F3EFECE9E6E3E0DDDAD7D4D1CECBC8C5C2BFBCB9B5B2AFACA9A6A3A09D9A97";
constant INIT_H_IBIA_22 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0C0C0C";
constant INIT_L_IBIA_22 : bit_vector(255 downto 0) := X"5754514E4B4845423F3C393633302D292623201D1A1714110E0B080502FFFCF9";
constant INIT_H_IBIA_23 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_IBIA_23 : bit_vector(255 downto 0) := X"B9B6B3B0ADAAA7A4A19D9A9794918E8B8885827F7C797673706D6A6763605D5A";
constant INIT_H_IBIA_24 : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_IBIA_24 : bit_vector(255 downto 0) := X"1B1815110E0B080502FFFCF9F6F3F0EDEAE7E4E1DEDBD7D4D1CECBC8C5C2BFBC";
constant INIT_H_IBIA_25 : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_IBIA_25 : bit_vector(255 downto 0) := X"7C797673706D6A6764615E5B5855524F4B4845423F3C393633302D2A2724211E";
constant INIT_H_IBIA_26 : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_IBIA_26 : bit_vector(255 downto 0) := X"DEDBD8D5D2CFCCC9C6C2BFBCB9B6B3B0ADAAA7A4A19E9B9895928F8C8885827F";
constant INIT_H_IBIA_27 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_IBIA_27 : bit_vector(255 downto 0) := X"403D3A3633302D2A2724211E1B1815120F0C09060300FCF9F6F3F0EDEAE7E4E1";
constant INIT_H_IBIA_28 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_IBIA_28 : bit_vector(255 downto 0) := X"A19E9B9895928F8C898683807D7A7774706D6A6764615E5B5855524F4C494643";
constant INIT_H_IBIA_29 : bit_vector(255 downto 0) := X"10100F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_IBIA_29 : bit_vector(255 downto 0) := X"0300FDFAF7F4F1EEEBE8E4E1DEDBD8D5D2CFCCC9C6C3C0BDBAB7B4B1AEAAA7A4";
constant INIT_H_IBIA_2A : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_IBIA_2A : bit_vector(255 downto 0) := X"65625F5C5855524F4C494643403D3A3734312E2B2825221E1B1815120F0C0906";
constant INIT_H_IBIA_2B : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_IBIA_2B : bit_vector(255 downto 0) := X"C6C3C0BDBAB7B4B1AEABA8A5A29F9C9996928F8C898683807D7A7774716E6B68";
constant INIT_H_IBIA_2C : bit_vector(255 downto 0) := X"1111111111111111111111111111101010101010101010101010101010101010";
constant INIT_L_IBIA_2C : bit_vector(255 downto 0) := X"2825221F1C191613100D0A060300FDFAF7F4F1EEEBE8E5E2DFDCD9D6D3D0CCC9";
constant INIT_H_IBIA_2D : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_IBIA_2D : bit_vector(255 downto 0) := X"8A8784817E7A7774716E6B6865625F5C595653504D4A4744403D3A3734312E2B";
constant INIT_H_IBIA_2E : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_IBIA_2E : bit_vector(255 downto 0) := X"EBE8E5E2DFDCD9D6D3D0CDCAC7C4C1BEBBB8B4B1AEABA8A5A29F9C999693908D";
constant INIT_H_IBIA_2F : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212111111111111";
constant INIT_L_IBIA_2F : bit_vector(255 downto 0) := X"4D4A4744413E3B3835322F2C2825221F1C191613100D0A070401FEFBF8F5F2EE";
constant INIT_H_IBIA_30 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_IBIA_30 : bit_vector(255 downto 0) := X"AFACA9A6A3A09C999693908D8A8784817E7B7875726F6C6966625F5C59565350";
constant INIT_H_IBIA_31 : bit_vector(255 downto 0) := X"1313131313131212121212121212121212121212121212121212121212121212";
constant INIT_L_IBIA_31 : bit_vector(255 downto 0) := X"100D0A070401FEFBF8F5F2EFECE9E6E3E0DDDAD6D3D0CDCAC7C4C1BEBBB8B5B2";
constant INIT_H_IBIA_32 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_IBIA_32 : bit_vector(255 downto 0) := X"726F6C696663605D5A5754514D4A4744413E3B3835322F2C292623201D1A1714";
constant INIT_H_IBIA_33 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_IBIA_33 : bit_vector(255 downto 0) := X"D4D1CECBC8C5C1BEBBB8B5B2AFACA9A6A3A09D9A9794918E8B8784817E7B7875";
constant INIT_H_IBIA_34 : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141313131313131313131313131313";
constant INIT_L_IBIA_34 : bit_vector(255 downto 0) := X"35322F2C292623201D1A1714110E0B080502FFFBF8F5F2EFECE9E6E3E0DDDAD7";
constant INIT_H_IBIA_35 : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_IBIA_35 : bit_vector(255 downto 0) := X"9794918E8B8885827F7C7976736F6C696663605D5A5754514E4B4845423F3C39";
constant INIT_H_IBIA_36 : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_IBIA_36 : bit_vector(255 downto 0) := X"F9F6F3F0EDEAE7E3E0DDDAD7D4D1CECBC8C5C2BFBCB9B6B3B0ADA9A6A3A09D9A";
constant INIT_H_IBIA_37 : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151414";
constant INIT_L_IBIA_37 : bit_vector(255 downto 0) := X"5B5754514E4B4845423F3C393633302D2A2724211D1A1714110E0B080502FFFC";
constant INIT_H_IBIA_38 : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_IBIA_38 : bit_vector(255 downto 0) := X"BCB9B6B3B0ADAAA7A4A19E9B9895918E8B8885827F7C797673706D6A6764615E";
constant INIT_H_IBIA_39 : bit_vector(255 downto 0) := X"1616161616161616161615151515151515151515151515151515151515151515";
constant INIT_L_IBIA_39 : bit_vector(255 downto 0) := X"1E1B1815120F0C090502FFFCF9F6F3F0EDEAE7E4E1DEDBD8D5D2CFCBC8C5C2BF";
constant INIT_H_IBIA_3A : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161616161616";
constant INIT_L_IBIA_3A : bit_vector(255 downto 0) := X"807D797673706D6A6764615E5B5855524F4C4946433F3C393633302D2A272421";
constant INIT_H_IBIA_3B : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161616161616";
constant INIT_L_IBIA_3B : bit_vector(255 downto 0) := X"E1DEDBD8D5D2CFCCC9C6C3C0BDBAB7B3B0ADAAA7A4A19E9B9895928F8C898683";
constant INIT_H_IBIA_3C : bit_vector(255 downto 0) := X"1717171717171717171717171717171717171717171717161616161616161616";
constant INIT_L_IBIA_3C : bit_vector(255 downto 0) := X"43403D3A3734312E2B2724211E1B1815120F0C09060300FDFAF7F4F1EDEAE7E4";
constant INIT_H_IBIA_3D : bit_vector(255 downto 0) := X"1717171717171717171717171717171717171717171717171717171717171717";
constant INIT_L_IBIA_3D : bit_vector(255 downto 0) := X"A5A29F9B9895928F8C898683807D7A7774716E6B6865615E5B5855524F4C4946";
constant INIT_H_IBIA_3E : bit_vector(255 downto 0) := X"1818181717171717171717171717171717171717171717171717171717171717";
constant INIT_L_IBIA_3E : bit_vector(255 downto 0) := X"060300FDFAF7F4F1EEEBE8E5E2DFDCD9D5D2CFCCC9C6C3C0BDBAB7B4B1AEABA8";
constant INIT_H_IBIA_3F : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_IBIA_3F : bit_vector(255 downto 0) := X"6865625F5C595653504C494643403D3A3734312E2B2825221F1C1916120F0C09";
constant INIT_H_IBIA_40 : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_IBIA_40 : bit_vector(255 downto 0) := X"CAC7C4C0BDBAB7B4B1AEABA8A5A29F9C999693908D8A8683807D7A7774716E6B";
constant INIT_H_IBIA_41 : bit_vector(255 downto 0) := X"1919191919191919191919191919191818181818181818181818181818181818";
constant INIT_L_IBIA_41 : bit_vector(255 downto 0) := X"2B2825221F1C191613100D0A070401FEFAF7F4F1EEEBE8E5E2DFDCD9D6D3D0CD";
constant INIT_H_IBIA_42 : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_IBIA_42 : bit_vector(255 downto 0) := X"8D8A8784817E7B7875726E6B6865625F5C595653504D4A4744413E3B3834312E";
constant INIT_H_IBIA_43 : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_IBIA_43 : bit_vector(255 downto 0) := X"EFECE9E6E2DFDCD9D6D3D0CDCAC7C4C1BEBBB8B5B2AFACA8A5A29F9C99969390";
constant INIT_H_IBIA_44 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1919191919";
constant INIT_L_IBIA_44 : bit_vector(255 downto 0) := X"504D4A4744413E3B3835322F2C292623201C191613100D0A070401FEFBF8F5F2";
constant INIT_H_IBIA_45 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_IBIA_45 : bit_vector(255 downto 0) := X"B2AFACA9A6A3A09D9A9794908D8A8784817E7B7875726F6C696663605D5A5653";
constant INIT_H_IBIA_46 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_IBIA_46 : bit_vector(255 downto 0) := X"14110E0B080401FEFBF8F5F2EFECE9E6E3E0DDDAD7D4D1CECAC7C4C1BEBBB8B5";
constant INIT_H_IBIA_47 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_IBIA_47 : bit_vector(255 downto 0) := X"75726F6C696663605D5A5754514E4B4845423E3B3835322F2C292623201D1A17";
constant INIT_H_IBIA_48 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_IBIA_48 : bit_vector(255 downto 0) := X"D7D4D1CECBC8C5C2BFBCB9B6B2AFACA9A6A3A09D9A9794918E8B8885827F7C78";
constant INIT_H_IBIA_49 : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_IBIA_49 : bit_vector(255 downto 0) := X"393633302D2A2623201D1A1714110E0B080502FFFCF9F6F3F0ECE9E6E3E0DDDA";
constant INIT_H_IBIA_4A : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_IBIA_4A : bit_vector(255 downto 0) := X"9A9794918E8B8885827F7C797673706D6A6764605D5A5754514E4B4845423F3C";
constant INIT_H_IBIA_4B : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_IBIA_4B : bit_vector(255 downto 0) := X"FCF9F6F3F0EDEAE7E4E1DEDBD7D4D1CECBC8C5C2BFBCB9B6B3B0ADAAA7A4A19E";
constant INIT_H_IBIA_4C : bit_vector(255 downto 0) := X"1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1C";
constant INIT_L_IBIA_4C : bit_vector(255 downto 0) := X"5E5B5855524F4B4845423F3C393633302D2A2724211E1B1815110E0B080502FF";
constant INIT_H_IBIA_4D : bit_vector(255 downto 0) := X"1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D";
constant INIT_L_IBIA_4D : bit_vector(255 downto 0) := X"BFBCB9B6B3B0ADAAA7A4A19E9B9895928F8C8985827F7C797673706D6A676461";
constant INIT_H_IBIA_4E : bit_vector(255 downto 0) := X"1E1E1E1E1E1E1E1E1E1E1E1E1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D";
constant INIT_L_IBIA_4E : bit_vector(255 downto 0) := X"211E1B1815120F0C09060300FDF9F6F3F0EDEAE7E4E1DEDBD8D5D2CFCCC9C6C3";
constant INIT_H_IBIA_4F : bit_vector(255 downto 0) := X"1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E";
constant INIT_L_IBIA_4F : bit_vector(255 downto 0) := X"83807D7A7774716D6A6764615E5B5855524F4C494643403D3A3733302D2A2724";
constant INIT_H_IBIA_50 : bit_vector(255 downto 0) := X"1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E";
constant INIT_L_IBIA_50 : bit_vector(255 downto 0) := X"E5E1DEDBD8D5D2CFCCC9C6C3C0BDBAB7B4B1AEABA7A4A19E9B9895928F8C8986";
constant INIT_H_IBIA_51 : bit_vector(255 downto 0) := X"1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1E1E1E1E1E1E1E1E";
constant INIT_L_IBIA_51 : bit_vector(255 downto 0) := X"4643403D3A3734312E2B2825221F1B1815120F0C09060300FDFAF7F4F1EEEBE8";
constant INIT_H_IBIA_52 : bit_vector(255 downto 0) := X"1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F";
constant INIT_L_IBIA_52 : bit_vector(255 downto 0) := X"A8A5A29F9C9996938F8C898683807D7A7774716E6B6865625F5C5955524F4C49";
constant INIT_H_IBIA_53 : bit_vector(255 downto 0) := X"202020201F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F";
constant INIT_L_IBIA_53 : bit_vector(255 downto 0) := X"0A070300FDFAF7F4F1EEEBE8E5E2DFDCD9D6D3D0CDC9C6C3C0BDBAB7B4B1AEAB";
constant INIT_H_IBIA_54 : bit_vector(255 downto 0) := X"2020202020202020202020202020202020202020202020202020202020202020";
constant INIT_L_IBIA_54 : bit_vector(255 downto 0) := X"6B6865625F5C595653504D4A4744413D3A3734312E2B2825221F1C191613100D";
constant INIT_H_IBIA_55 : bit_vector(255 downto 0) := X"2020202020202020202020202020202020202020202020202020202020202020";
constant INIT_L_IBIA_55 : bit_vector(255 downto 0) := X"CDCAC7C4C1BEBBB8B5B1AEABA8A5A29F9C999693908D8A8784817E7B7774716E";
constant INIT_H_IBIA_56 : bit_vector(255 downto 0) := X"2121212121212121212121212121212120202020202020202020202020202020";
constant INIT_L_IBIA_56 : bit_vector(255 downto 0) := X"2F2C2925221F1C191613100D0A070401FEFBF8F5F2EFEBE8E5E2DFDCD9D6D3D0";
constant INIT_H_IBIA_57 : bit_vector(255 downto 0) := X"2121212121212121212121212121212121212121212121212121212121212121";
constant INIT_L_IBIA_57 : bit_vector(255 downto 0) := X"908D8A8784817E7B7875726F6C6966635F5C595653504D4A4744413E3B383532";
constant INIT_H_IBIA_58 : bit_vector(255 downto 0) := X"2121212121212121212121212121212121212121212121212121212121212121";
constant INIT_L_IBIA_58 : bit_vector(255 downto 0) := X"F2EFECE9E6E3E0DDDAD6D3D0CDCAC7C4C1BEBBB8B5B2AFACA9A6A3A09C999693";
constant INIT_H_IBIA_59 : bit_vector(255 downto 0) := X"2222222222222222222222222222222222222222222222222222222221212121";
constant INIT_L_IBIA_59 : bit_vector(255 downto 0) := X"54514E4A4744413E3B3835322F2C292623201D1A1714100D0A070401FEFBF8F5";
constant INIT_H_IBIA_5A : bit_vector(255 downto 0) := X"2222222222222222222222222222222222222222222222222222222222222222";
constant INIT_L_IBIA_5A : bit_vector(255 downto 0) := X"B5B2AFACA9A6A3A09D9A9794918E8B8884817E7B7875726F6C696663605D5A57";
constant INIT_H_IBIA_5B : bit_vector(255 downto 0) := X"2323232323232323222222222222222222222222222222222222222222222222";
constant INIT_L_IBIA_5B : bit_vector(255 downto 0) := X"1714110E0B080502FFFCF8F5F2EFECE9E6E3E0DDDAD7D4D1CECBC8C5C2BEBBB8";
constant INIT_H_IBIA_5C : bit_vector(255 downto 0) := X"2323232323232323232323232323232323232323232323232323232323232323";
constant INIT_L_IBIA_5C : bit_vector(255 downto 0) := X"797673706C696663605D5A5754514E4B4845423F3C3936322F2C292623201D1A";
constant INIT_H_IBIA_5D : bit_vector(255 downto 0) := X"2323232323232323232323232323232323232323232323232323232323232323";
constant INIT_L_IBIA_5D : bit_vector(255 downto 0) := X"DAD7D4D1CECBC8C5C2BFBCB9B6B3B0ADAAA6A3A09D9A9794918E8B8885827F7C";
constant INIT_H_IBIA_5E : bit_vector(255 downto 0) := X"2424242424242424242424242424242424242424232323232323232323232323";
constant INIT_L_IBIA_5E : bit_vector(255 downto 0) := X"3C393633302D2A2724211E1A1714110E0B080502FFFCF9F6F3F0EDEAE7E4E0DD";
constant INIT_H_IBIA_5F : bit_vector(255 downto 0) := X"2424242424242424242424242424242424242424242424242424242424242424";
constant INIT_L_IBIA_5F : bit_vector(255 downto 0) := X"9E9B9895928E8B8885827F7C797673706D6A6764615E5B5854514E4B4845423F";
constant INIT_H_IBIA_60 : bit_vector(255 downto 0) := X"2424242424242424242424242424242424242424242424242424242424242424";
constant INIT_L_IBIA_60 : bit_vector(255 downto 0) := X"FFFCF9F6F3F0EDEAE7E4E1DEDBD8D5D2CFCCC8C5C2BFBCB9B6B3B0ADAAA7A4A1";
constant INIT_H_IBIA_61 : bit_vector(255 downto 0) := X"2525252525252525252525252525252525252525252525252525252525252525";
constant INIT_L_IBIA_61 : bit_vector(255 downto 0) := X"615E5B5855524F4C494643403C393633302D2A2724211E1B1815120F0C090602";
constant INIT_H_IBIA_62 : bit_vector(255 downto 0) := X"2525252525252525252525252525252525252525252525252525252525252525";
constant INIT_L_IBIA_62 : bit_vector(255 downto 0) := X"C3C0BDBAB7B4B0ADAAA7A4A19E9B9895928F8C898683807D7A7673706D6A6764";
constant INIT_H_IBIA_63 : bit_vector(255 downto 0) := X"2626262626262626262626262625252525252525252525252525252525252525";
constant INIT_L_IBIA_63 : bit_vector(255 downto 0) := X"24211E1B1815120F0C09060300FDFAF7F4F1EEEAE7E4E1DEDBD8D5D2CFCCC9C6";
constant INIT_H_IBIA_64 : bit_vector(255 downto 0) := X"2626262626262626262626262626262626262626262626262626262626262626";
constant INIT_L_IBIA_64 : bit_vector(255 downto 0) := X"8683807D7A7774716E6B6865615E5B5855524F4C494643403D3A3734312E2B28";
constant INIT_H_IBIA_65 : bit_vector(255 downto 0) := X"2626262626262626262626262626262626262626262626262626262626262626";
constant INIT_L_IBIA_65 : bit_vector(255 downto 0) := X"E8E5E2DFDCD9D5D2CFCCC9C6C3C0BDBAB7B4B1AEABA8A5A29F9B9895928F8C89";
constant INIT_H_IBIA_66 : bit_vector(255 downto 0) := X"2727272727272727272727272727272727272727272727272726262626262626";
constant INIT_L_IBIA_66 : bit_vector(255 downto 0) := X"494643403D3A3734312E2B2825221F1C1916130F0C09060300FDFAF7F4F1EEEB";
constant INIT_H_IBIA_67 : bit_vector(255 downto 0) := X"2727272727272727272727272727272727272727272727272727272727272727";
constant INIT_L_IBIA_67 : bit_vector(255 downto 0) := X"ABA8A5A29F9C999693908D8A8783807D7A7774716E6B6865625F5C595653504D";
constant INIT_H_IBIA_68 : bit_vector(255 downto 0) := X"2828282828272727272727272727272727272727272727272727272727272727";
constant INIT_L_IBIA_68 : bit_vector(255 downto 0) := X"0D0A070401FEFBF7F4F1EEEBE8E5E2DFDCD9D6D3D0CDCAC7C4C1BDBAB7B4B1AE";
constant INIT_H_IBIA_69 : bit_vector(255 downto 0) := X"2828282828282828282828282828282828282828282828282828282828282828";
constant INIT_L_IBIA_69 : bit_vector(255 downto 0) := X"6F6B6865625F5C595653504D4A4744413E3B3835312E2B2825221F1C19161310";
constant INIT_H_IBIA_6A : bit_vector(255 downto 0) := X"2828282828282828282828282828282828282828282828282828282828282828";
constant INIT_L_IBIA_6A : bit_vector(255 downto 0) := X"D0CDCAC7C4C1BEBBB8B5B2AFACA9A5A29F9C999693908D8A8784817E7B787572";
constant INIT_H_IBIA_6B : bit_vector(255 downto 0) := X"2929292929292929292929292929292929282828282828282828282828282828";
constant INIT_L_IBIA_6B : bit_vector(255 downto 0) := X"322F2C292623201D191613100D0A070401FEFBF8F5F2EFECE9E6E3DFDCD9D6D3";
constant INIT_H_IBIA_6C : bit_vector(255 downto 0) := X"2929292929292929292929292929292929292929292929292929292929292929";
constant INIT_L_IBIA_6C : bit_vector(255 downto 0) := X"94918D8A8784817E7B7875726F6C696663605D5A5753504D4A4744413E3B3835";
constant INIT_H_IBIA_6D : bit_vector(255 downto 0) := X"2929292929292929292929292929292929292929292929292929292929292929";
constant INIT_L_IBIA_6D : bit_vector(255 downto 0) := X"F5F2EFECE9E6E3E0DDDAD7D4D1CECBC7C4C1BEBBB8B5B2AFACA9A6A3A09D9A97";
constant INIT_H_IBIA_6E : bit_vector(255 downto 0) := X"2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A292929";
constant INIT_L_IBIA_6E : bit_vector(255 downto 0) := X"5754514E4B4845423F3B3835322F2C292623201D1A1714110E0B080501FEFBF8";
constant INIT_H_IBIA_6F : bit_vector(255 downto 0) := X"2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A";
constant INIT_L_IBIA_6F : bit_vector(255 downto 0) := X"B9B6B3AFACA9A6A3A09D9A9794918E8B8885827F7C7975726F6C696663605D5A";
constant INIT_H_IBIA_70 : bit_vector(255 downto 0) := X"2B2B2B2B2B2B2B2B2B2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A";
constant INIT_L_IBIA_70 : bit_vector(255 downto 0) := X"1A1714110E0B080502FFFCF9F6F3F0EDE9E6E3E0DDDAD7D4D1CECBC8C5C2BFBC";
constant INIT_H_IBIA_71 : bit_vector(255 downto 0) := X"2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B";
constant INIT_L_IBIA_71 : bit_vector(255 downto 0) := X"7C797673706D6A6764605D5A5754514E4B4845423F3C393633302D2A2623201D";
constant INIT_H_IBIA_72 : bit_vector(255 downto 0) := X"2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B";
constant INIT_L_IBIA_72 : bit_vector(255 downto 0) := X"DEDBD8D4D1CECBC8C5C2BFBCB9B6B3B0ADAAA7A4A19E9A9794918E8B8885827F";
constant INIT_H_IBIA_73 : bit_vector(255 downto 0) := X"2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2B2B2B2B2B2B2B2B2B2B2B";
constant INIT_L_IBIA_73 : bit_vector(255 downto 0) := X"3F3C393633302D2A2724211E1B1815120E0B080502FFFCF9F6F3F0EDEAE7E4E1";
constant INIT_H_IBIA_74 : bit_vector(255 downto 0) := X"2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C";
constant INIT_L_IBIA_74 : bit_vector(255 downto 0) := X"A19E9B9895928F8C8986827F7C797673706D6A6764615E5B5855524F4C484542";
constant INIT_H_IBIA_75 : bit_vector(255 downto 0) := X"2D2D2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C";
constant INIT_L_IBIA_75 : bit_vector(255 downto 0) := X"0300FDFAF6F3F0EDEAE7E4E1DEDBD8D5D2CFCCC9C6C3C0BCB9B6B3B0ADAAA7A4";
constant INIT_H_IBIA_76 : bit_vector(255 downto 0) := X"2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D";
constant INIT_L_IBIA_76 : bit_vector(255 downto 0) := X"64615E5B5855524F4C494643403D3A3734302D2A2724211E1B1815120F0C0906";
constant INIT_H_IBIA_77 : bit_vector(255 downto 0) := X"2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D";
constant INIT_L_IBIA_77 : bit_vector(255 downto 0) := X"C6C3C0BDBAB7B4B1AEABA8A4A19E9B9895928F8C898683807D7A7774716E6A67";
constant INIT_H_IBIA_78 : bit_vector(255 downto 0) := X"2E2E2E2E2E2E2E2E2E2E2E2E2E2E2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D";
constant INIT_L_IBIA_78 : bit_vector(255 downto 0) := X"2825221F1C1815120F0C09060300FDFAF7F4F1EEEBE8E5E2DEDBD8D5D2CFCCC9";
constant INIT_H_IBIA_79 : bit_vector(255 downto 0) := X"2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E";
constant INIT_L_IBIA_79 : bit_vector(255 downto 0) := X"898683807D7A7774716E6B6865625F5C5956524F4C494643403D3A3734312E2B";
constant INIT_H_IBIA_7A : bit_vector(255 downto 0) := X"2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E";
constant INIT_L_IBIA_7A : bit_vector(255 downto 0) := X"EBE8E5E2DFDCD9D6D3D0CDCAC6C3C0BDBAB7B4B1AEABA8A5A29F9C999693908C";
constant INIT_H_IBIA_7B : bit_vector(255 downto 0) := X"2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2E2E2E2E2E2E";
constant INIT_L_IBIA_7B : bit_vector(255 downto 0) := X"4D4A4744413E3A3734312E2B2825221F1C191613100D0A070400FDFAF7F4F1EE";
constant INIT_H_IBIA_7C : bit_vector(255 downto 0) := X"2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F";
constant INIT_L_IBIA_7C : bit_vector(255 downto 0) := X"AEABA8A5A29F9C999693908D8A8784817E7B7874716E6B6865625F5C59565350";
constant INIT_H_IBIA_7D : bit_vector(255 downto 0) := X"3030303030302F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F";
constant INIT_L_IBIA_7D : bit_vector(255 downto 0) := X"100D0A070401FEFBF8F5F2EFEBE8E5E2DFDCD9D6D3D0CDCAC7C4C1BEBBB8B5B2";
constant INIT_H_IBIA_7E : bit_vector(255 downto 0) := X"3030303030303030303030303030303030303030303030303030303030303030";
constant INIT_L_IBIA_7E : bit_vector(255 downto 0) := X"726F6C6966635F5C595653504D4A4744413E3B3835322F2C2925221F1C191613";
constant INIT_H_IBIA_7F : bit_vector(255 downto 0) := X"3030303030303030303030303030303030303030303030303030303030303030";
constant INIT_L_IBIA_7F : bit_vector(255 downto 0) := X"D3D0CDCAC7C4C1BEBBB8B5B2AFACA9A6A3A09D999693908D8A8784817E7B7875";
constant INIT_H_AVIN_00 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_AVIN_00 : bit_vector(255 downto 0) := X"38363533312F2D2B2A28262422201F1D1B1917151412100E0C0A090705030100";
constant INIT_H_AVIN_01 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_AVIN_01 : bit_vector(255 downto 0) := X"73716F6D6C6A68666462615F5D5B5957565452504E4C4B4947454341403E3C3A";
constant INIT_H_AVIN_02 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_AVIN_02 : bit_vector(255 downto 0) := X"ADACAAA8A6A4A3A19F9D9B9998969492908E8D8B8987858382807E7C7A787775";
constant INIT_H_AVIN_03 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_AVIN_03 : bit_vector(255 downto 0) := X"E8E6E4E3E1DFDDDBD9D8D6D4D2D0CECDCBC9C7C5C3C2C0BEBCBAB8B7B5B3B1AF";
constant INIT_H_AVIN_04 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101000000000000000000000000";
constant INIT_L_AVIN_04 : bit_vector(255 downto 0) := X"23211F1D1B1A18161412100F0D0B090705040200FEFCFAF9F7F5F3F1EFEEECEA";
constant INIT_H_AVIN_05 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_AVIN_05 : bit_vector(255 downto 0) := X"5D5B5A58565452504F4D4B4947464442403E3C3B3937353331302E2C2A282625";
constant INIT_H_AVIN_06 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_AVIN_06 : bit_vector(255 downto 0) := X"98969492918F8D8B8987868482807E7C7B7977757371706E6C6A68666563615F";
constant INIT_H_AVIN_07 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_AVIN_07 : bit_vector(255 downto 0) := X"D3D1CFCDCBC9C8C6C4C2C0BEBDBBB9B7B5B3B2B0AEACAAA8A7A5A3A19F9D9C9A";
constant INIT_H_AVIN_08 : bit_vector(255 downto 0) := X"0202020202020202010101010101010101010101010101010101010101010101";
constant INIT_L_AVIN_08 : bit_vector(255 downto 0) := X"0D0B090806040200FEFDFBF9F7F5F4F2F0EEECEAE9E7E5E3E1DFDEDCDAD8D6D4";
constant INIT_H_AVIN_09 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_AVIN_09 : bit_vector(255 downto 0) := X"48464442403F3D3B3937353432302E2C2A29272523211F1E1C1A18161413110F";
constant INIT_H_AVIN_0A : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_AVIN_0A : bit_vector(255 downto 0) := X"82817F7D7B7977767472706E6C6B6967656361605E5C5A58565553514F4D4B4A";
constant INIT_H_AVIN_0B : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_AVIN_0B : bit_vector(255 downto 0) := X"BDBBB9B7B6B4B2B0AEACABA9A7A5A3A1A09E9C9A98979593918F8D8C8A888684";
constant INIT_H_AVIN_0C : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_AVIN_0C : bit_vector(255 downto 0) := X"F8F6F4F2F0EEEDEBE9E7E5E3E2E0DEDCDAD8D7D5D3D1CFCDCCCAC8C6C4C2C1BF";
constant INIT_H_AVIN_0D : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030302020202";
constant INIT_L_AVIN_0D : bit_vector(255 downto 0) := X"32302F2D2B2927252422201E1C1A19171513110F0E0C0A0806040301FFFDFBF9";
constant INIT_H_AVIN_0E : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_AVIN_0E : bit_vector(255 downto 0) := X"6D6B6967656462605E5C5A59575553514F4E4C4A48464443413F3D3B3A383634";
constant INIT_H_AVIN_0F : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_AVIN_0F : bit_vector(255 downto 0) := X"A7A6A4A2A09E9C9B9997959391908E8C8A88868583817F7D7B7A78767472706F";
constant INIT_H_AVIN_10 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_AVIN_10 : bit_vector(255 downto 0) := X"E2E0DEDDDBD9D7D5D3D2D0CECCCAC8C7C5C3C1BFBDBCBAB8B6B4B2B1AFADABA9";
constant INIT_H_AVIN_11 : bit_vector(255 downto 0) := X"0404040404040404040404040404040403030303030303030303030303030303";
constant INIT_L_AVIN_11 : bit_vector(255 downto 0) := X"1D1B1917151312100E0C0A0807050301FFFDFCFAF8F6F4F2F1EFEDEBE9E8E6E4";
constant INIT_H_AVIN_12 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_AVIN_12 : bit_vector(255 downto 0) := X"57555452504E4C4A49474543413F3E3C3A38363433312F2D2B2928262422201E";
constant INIT_H_AVIN_13 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_AVIN_13 : bit_vector(255 downto 0) := X"92908E8C8B8987858381807E7C7A78767573716F6D6B6A68666462605F5D5B59";
constant INIT_H_AVIN_14 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_AVIN_14 : bit_vector(255 downto 0) := X"CCCBC9C7C5C3C1C0BEBCBAB8B6B5B3B1AFADABAAA8A6A4A2A09F9D9B99979594";
constant INIT_H_AVIN_15 : bit_vector(255 downto 0) := X"0505050505040404040404040404040404040404040404040404040404040404";
constant INIT_L_AVIN_15 : bit_vector(255 downto 0) := X"0705030200FEFCFAF8F7F5F3F1EFEDECEAE8E6E4E2E1DFDDDBD9D7D6D4D2D0CE";
constant INIT_H_AVIN_16 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_AVIN_16 : bit_vector(255 downto 0) := X"42403E3C3A38373533312F2E2C2A28262423211F1D1B1918161412100E0D0B09";
constant INIT_H_AVIN_17 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_AVIN_17 : bit_vector(255 downto 0) := X"7C7A79777573716F6E6C6A68666463615F5D5B5958565452504E4D4B49474543";
constant INIT_H_AVIN_18 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_AVIN_18 : bit_vector(255 downto 0) := X"B7B5B3B1B0AEACAAA8A6A5A3A19F9D9B9A98969492908F8D8B8987858482807E";
constant INIT_H_AVIN_19 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_AVIN_19 : bit_vector(255 downto 0) := X"F1F0EEECEAE8E6E5E3E1DFDDDCDAD8D6D4D2D1CFCDCBC9C7C6C4C2C0BEBCBBB9";
constant INIT_H_AVIN_1A : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060605050505050505";
constant INIT_L_AVIN_1A : bit_vector(255 downto 0) := X"2C2A28272523211F1D1C1A18161412110F0D0B090706040200FEFCFBF9F7F5F3";
constant INIT_H_AVIN_1B : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_AVIN_1B : bit_vector(255 downto 0) := X"676563615F5E5C5A58565453514F4D4B4948464442403E3D3B3937353332302E";
constant INIT_H_AVIN_1C : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_AVIN_1C : bit_vector(255 downto 0) := X"A19F9E9C9A98969493918F8D8B8988868482807F7D7B7977757472706E6C6A69";
constant INIT_H_AVIN_1D : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_AVIN_1D : bit_vector(255 downto 0) := X"DCDAD8D6D5D3D1CFCDCBCAC8C6C4C2C0BFBDBBB9B7B5B4B2B0AEACAAA9A7A5A3";
constant INIT_H_AVIN_1E : bit_vector(255 downto 0) := X"0707070707070707070707070706060606060606060606060606060606060606";
constant INIT_L_AVIN_1E : bit_vector(255 downto 0) := X"171513110F0D0C0A0806040201FFFDFBF9F7F6F4F2F0EEECEBE9E7E5E3E1E0DE";
constant INIT_H_AVIN_1F : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_AVIN_1F : bit_vector(255 downto 0) := X"514F4D4C4A48464442413F3D3B3937363432302E2C2B2927252322201E1C1A18";
constant INIT_H_AVIN_20 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_AVIN_20 : bit_vector(255 downto 0) := X"8C8A88868483817F7D7B7978767472706E6D6B6967656362605E5C5A58575553";
constant INIT_H_AVIN_21 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_AVIN_21 : bit_vector(255 downto 0) := X"C6C5C3C1BFBDBBBAB8B6B4B2B0AFADABA9A7A5A4A2A09E9C9A99979593918F8E";
constant INIT_H_AVIN_22 : bit_vector(255 downto 0) := X"0807070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_AVIN_22 : bit_vector(255 downto 0) := X"01FFFDFBFAF8F6F4F2F0EFEDEBE9E7E5E4E2E0DEDCDAD9D7D5D3D1D0CECCCAC8";
constant INIT_H_AVIN_23 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_AVIN_23 : bit_vector(255 downto 0) := X"3C3A38363432312F2D2B2927262422201E1C1B1917151311100E0C0A08060503";
constant INIT_H_AVIN_24 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_AVIN_24 : bit_vector(255 downto 0) := X"767473716F6D6B6968666462605E5D5B5957555352504E4C4A48474543413F3D";
constant INIT_H_AVIN_25 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_AVIN_25 : bit_vector(255 downto 0) := X"B1AFADABA9A8A6A4A2A09E9D9B9997959392908E8C8A88878583817F7D7C7A78";
constant INIT_H_AVIN_26 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_AVIN_26 : bit_vector(255 downto 0) := X"EBEAE8E6E4E2E0DFDDDBD9D7D5D4D2D0CECCCAC9C7C5C3C1BFBEBCBAB8B6B4B3";
constant INIT_H_AVIN_27 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090908080808080808080808";
constant INIT_L_AVIN_27 : bit_vector(255 downto 0) := X"262422201F1D1B1917161412100E0C0B090705030100FEFCFAF8F6F5F3F1EFED";
constant INIT_H_AVIN_28 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_AVIN_28 : bit_vector(255 downto 0) := X"615F5D5B5957565452504E4C4B4947454341403E3C3A38363533312F2D2B2A28";
constant INIT_H_AVIN_29 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_AVIN_29 : bit_vector(255 downto 0) := X"9B9998969492908E8D8B8987858382807E7C7A78777573716F6D6C6A68666462";
constant INIT_H_AVIN_2A : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_AVIN_2A : bit_vector(255 downto 0) := X"D6D4D2D0CECDCBC9C7C5C4C2C0BEBCBAB9B7B5B3B1AFAEACAAA8A6A4A3A19F9D";
constant INIT_H_AVIN_2B : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A09090909090909090909090909090909090909090909";
constant INIT_L_AVIN_2B : bit_vector(255 downto 0) := X"100F0D0B090705040200FEFCFAF9F7F5F3F1EFEEECEAE8E6E4E3E1DFDDDBD9D8";
constant INIT_H_AVIN_2C : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_AVIN_2C : bit_vector(255 downto 0) := X"4B4947464442403E3C3B3937353331302E2C2A28262523211F1D1B1A18161412";
constant INIT_H_AVIN_2D : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_AVIN_2D : bit_vector(255 downto 0) := X"868482807E7C7B7977757371706E6C6A68676563615F5D5C5A58565452514F4D";
constant INIT_H_AVIN_2E : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_AVIN_2E : bit_vector(255 downto 0) := X"C0BEBDBBB9B7B5B3B2B0AEACAAA8A7A5A3A19F9D9C9A98969492918F8D8B8987";
constant INIT_H_AVIN_2F : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_AVIN_2F : bit_vector(255 downto 0) := X"FBF9F7F5F4F2F0EEECEAE9E7E5E3E1DFDEDCDAD8D6D4D3D1CFCDCBC9C8C6C4C2";
constant INIT_H_AVIN_30 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0A0A";
constant INIT_L_AVIN_30 : bit_vector(255 downto 0) := X"353432302E2C2A29272523211F1E1C1A18161413110F0D0B0A0806040200FFFD";
constant INIT_H_AVIN_31 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_AVIN_31 : bit_vector(255 downto 0) := X"706E6C6B6967656361605E5C5A58565553514F4D4B4A48464442403F3D3B3937";
constant INIT_H_AVIN_32 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_AVIN_32 : bit_vector(255 downto 0) := X"ABA9A7A5A3A2A09E9C9A98979593918F8D8C8A88868482817F7D7B7977767472";
constant INIT_H_AVIN_33 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_AVIN_33 : bit_vector(255 downto 0) := X"E5E3E2E0DEDCDAD8D7D5D3D1CFCDCCCAC8C6C4C2C1BFBDBBB9B8B6B4B2B0AEAD";
constant INIT_H_AVIN_34 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_AVIN_34 : bit_vector(255 downto 0) := X"201E1C1A19171513110F0E0C0A0806040301FFFDFBF9F8F6F4F2F0EEEDEBE9E7";
constant INIT_H_AVIN_35 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_AVIN_35 : bit_vector(255 downto 0) := X"5B5957555351504E4C4A48464543413F3D3B3A38363432302F2D2B2927252422";
constant INIT_H_AVIN_36 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_AVIN_36 : bit_vector(255 downto 0) := X"959391908E8C8A88868583817F7D7B7A78767472706F6D6B6967656462605E5C";
constant INIT_H_AVIN_37 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_AVIN_37 : bit_vector(255 downto 0) := X"D0CECCCAC8C7C5C3C1BFBDBCBAB8B6B4B2B1AFADABA9A7A6A4A2A09E9C9B9997";
constant INIT_H_AVIN_38 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_AVIN_38 : bit_vector(255 downto 0) := X"0A0807050301FFFEFCFAF8F6F4F3F1EFEDEBE9E8E6E4E2E0DEDDDBD9D7D5D3D2";
constant INIT_H_AVIN_39 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_AVIN_39 : bit_vector(255 downto 0) := X"4543413F3E3C3A38363433312F2D2B2928262422201E1D1B1917151312100E0C";
constant INIT_H_AVIN_3A : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_AVIN_3A : bit_vector(255 downto 0) := X"807E7C7A78767573716F6D6B6A68666462605F5D5B5957555452504E4C4A4947";
constant INIT_H_AVIN_3B : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_AVIN_3B : bit_vector(255 downto 0) := X"BAB8B6B5B3B1AFADACAAA8A6A4A2A19F9D9B9997969492908E8C8B8987858381";
constant INIT_H_AVIN_3C : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_AVIN_3C : bit_vector(255 downto 0) := X"F5F3F1EFEDECEAE8E6E4E2E1DFDDDBD9D7D6D4D2D0CECCCBC9C7C5C3C1C0BEBC";
constant INIT_H_AVIN_3D : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0D0D0D0D0D";
constant INIT_L_AVIN_3D : bit_vector(255 downto 0) := X"2F2E2C2A28262423211F1D1B1918161412100E0D0B090705030200FEFCFAF8F7";
constant INIT_H_AVIN_3E : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_AVIN_3E : bit_vector(255 downto 0) := X"6A68666463615F5D5B5958565452504F4D4B4947454442403E3C3A3937353331";
constant INIT_H_AVIN_3F : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_AVIN_3F : bit_vector(255 downto 0) := X"A5A3A19F9D9B9A98969492908F8D8B8987858482807E7C7A79777573716F6E6C";
constant INIT_H_AVIN_40 : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_AVIN_40 : bit_vector(255 downto 0) := X"DFDDDCDAD8D6D4D2D1CFCDCBC9C7C6C4C2C0BEBCBBB9B7B5B3B1B0AEACAAA8A6";
constant INIT_H_AVIN_41 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_AVIN_41 : bit_vector(255 downto 0) := X"1A18161412110F0D0B090706040200FEFCFBF9F7F5F3F2F0EEECEAE8E7E5E3E1";
constant INIT_H_AVIN_42 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_AVIN_42 : bit_vector(255 downto 0) := X"5453514F4D4B4948464442403E3D3B3937353332302E2C2A28272523211F1D1C";
constant INIT_H_AVIN_43 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_AVIN_43 : bit_vector(255 downto 0) := X"8F8D8B8A88868482807F7D7B7977757472706E6C6A69676563615F5E5C5A5856";
constant INIT_H_AVIN_44 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_AVIN_44 : bit_vector(255 downto 0) := X"CAC8C6C4C2C0BFBDBBB9B7B5B4B2B0AEACAAA9A7A5A3A1A09E9C9A9896959391";
constant INIT_H_AVIN_45 : bit_vector(255 downto 0) := X"1010100F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_AVIN_45 : bit_vector(255 downto 0) := X"040201FFFDFBF9F7F6F4F2F0EEECEBE9E7E5E3E1E0DEDCDAD8D6D5D3D1CFCDCB";
constant INIT_H_AVIN_46 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_AVIN_46 : bit_vector(255 downto 0) := X"3F3D3B3938363432302E2D2B2927252322201E1C1A18171513110F0D0C0A0806";
constant INIT_H_AVIN_47 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_AVIN_47 : bit_vector(255 downto 0) := X"7978767472706E6D6B6967656362605E5C5A58575553514F4D4C4A4846444341";
constant INIT_H_AVIN_48 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_AVIN_48 : bit_vector(255 downto 0) := X"B4B2B0AFADABA9A7A5A4A2A09E9C9A99979593918F8E8C8A88868483817F7D7B";
constant INIT_H_AVIN_49 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_AVIN_49 : bit_vector(255 downto 0) := X"EFEDEBE9E7E6E4E2E0DEDCDBD9D7D5D3D1D0CECCCAC8C6C5C3C1BFBDBBBAB8B6";
constant INIT_H_AVIN_4A : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111101010101010101010";
constant INIT_L_AVIN_4A : bit_vector(255 downto 0) := X"2927262422201E1C1B1917151311100E0C0A0806050301FFFDFBFAF8F6F4F2F0";
constant INIT_H_AVIN_4B : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_AVIN_4B : bit_vector(255 downto 0) := X"6462605E5D5B5957555352504E4C4A48474543413F3D3C3A38363432312F2D2B";
constant INIT_H_AVIN_4C : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_AVIN_4C : bit_vector(255 downto 0) := X"9E9D9B9997959492908E8C8A89878583817F7E7C7A78767473716F6D6B696866";
constant INIT_H_AVIN_4D : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_AVIN_4D : bit_vector(255 downto 0) := X"D9D7D5D4D2D0CECCCAC9C7C5C3C1BFBEBCBAB8B6B4B3B1AFADABA9A8A6A4A2A0";
constant INIT_H_AVIN_4E : bit_vector(255 downto 0) := X"1212121212121212121212121111111111111111111111111111111111111111";
constant INIT_L_AVIN_4E : bit_vector(255 downto 0) := X"1412100E0C0B090705030100FEFCFAF8F6F5F3F1EFEDEBEAE8E6E4E2E0DFDDDB";
constant INIT_H_AVIN_4F : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_AVIN_4F : bit_vector(255 downto 0) := X"4E4C4B4947454341403E3C3A38373533312F2D2C2A28262422211F1D1B191716";
constant INIT_H_AVIN_50 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_AVIN_50 : bit_vector(255 downto 0) := X"8987858382807E7C7A78777573716F6D6C6A68666462615F5D5B595756545250";
constant INIT_H_AVIN_51 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_AVIN_51 : bit_vector(255 downto 0) := X"C4C2C0BEBCBAB9B7B5B3B1AFAEACAAA8A6A4A3A19F9D9B9998969492908E8D8B";
constant INIT_H_AVIN_52 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_AVIN_52 : bit_vector(255 downto 0) := X"FEFCFAF9F7F5F3F1EFEEECEAE8E6E4E3E1DFDDDBDAD8D6D4D2D0CFCDCBC9C7C5";
constant INIT_H_AVIN_53 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_AVIN_53 : bit_vector(255 downto 0) := X"3937353331302E2C2A28262523211F1D1B1A18161412100F0D0B090705040200";
constant INIT_H_AVIN_54 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_AVIN_54 : bit_vector(255 downto 0) := X"7372706E6C6A68676563615F5D5C5A58565452514F4D4B4947464442403E3C3B";
constant INIT_H_AVIN_55 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_AVIN_55 : bit_vector(255 downto 0) := X"AEACAAA8A7A5A3A19F9D9C9A98969492918F8D8B8988868482807E7D7B797775";
constant INIT_H_AVIN_56 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_AVIN_56 : bit_vector(255 downto 0) := X"E9E7E5E3E1DFDEDCDAD8D6D4D3D1CFCDCBC9C8C6C4C2C0BEBDBBB9B7B5B3B2B0";
constant INIT_H_AVIN_57 : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414131313131313131313131313";
constant INIT_L_AVIN_57 : bit_vector(255 downto 0) := X"2321201E1C1A18161513110F0D0B0A0806040200FFFDFBF9F7F5F4F2F0EEECEA";
constant INIT_H_AVIN_58 : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_AVIN_58 : bit_vector(255 downto 0) := X"5E5C5A58565553514F4D4B4A48464442403F3D3B3937353432302E2C2B292725";
constant INIT_H_AVIN_59 : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_AVIN_59 : bit_vector(255 downto 0) := X"98979593918F8D8C8A88868482817F7D7B7977767472706E6C6B696765636160";
constant INIT_H_AVIN_5A : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_AVIN_5A : bit_vector(255 downto 0) := X"D3D1CFCECCCAC8C6C4C3C1BFBDBBB9B8B6B4B2B0AEADABA9A7A5A3A2A09E9C9A";
constant INIT_H_AVIN_5B : bit_vector(255 downto 0) := X"1515151515151515141414141414141414141414141414141414141414141414";
constant INIT_L_AVIN_5B : bit_vector(255 downto 0) := X"0E0C0A0806040301FFFDFBF9F8F6F4F2F0EEEDEBE9E7E5E3E2E0DEDCDAD8D7D5";
constant INIT_H_AVIN_5C : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_AVIN_5C : bit_vector(255 downto 0) := X"48464543413F3D3B3A38363432302F2D2B2927252422201E1C1A19171513110F";
constant INIT_H_AVIN_5D : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_AVIN_5D : bit_vector(255 downto 0) := X"83817F7D7C7A78767472716F6D6B6967666462605E5C5B5957555351504E4C4A";
constant INIT_H_AVIN_5E : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_AVIN_5E : bit_vector(255 downto 0) := X"BDBCBAB8B6B4B2B1AFADABA9A7A6A4A2A09E9C9B9997959391908E8C8A888685";
constant INIT_H_AVIN_5F : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_AVIN_5F : bit_vector(255 downto 0) := X"F8F6F4F3F1EFEDEBE9E8E6E4E2E0DEDDDBD9D7D5D3D2D0CECCCAC8C7C5C3C1BF";
constant INIT_H_AVIN_60 : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161615151515";
constant INIT_L_AVIN_60 : bit_vector(255 downto 0) := X"33312F2D2B2928262422201F1D1B1917151412100E0C0A0907050301FFFEFCFA";
constant INIT_H_AVIN_61 : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161616161616";
constant INIT_L_AVIN_61 : bit_vector(255 downto 0) := X"6D6B6A68666462605F5D5B5957555452504E4C4A49474543413F3E3C3A383634";
constant INIT_H_AVIN_62 : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161616161616";
constant INIT_L_AVIN_62 : bit_vector(255 downto 0) := X"A8A6A4A2A19F9D9B9997969492908E8C8B8987858381807E7C7A78767573716F";
constant INIT_H_AVIN_63 : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161616161616";
constant INIT_L_AVIN_63 : bit_vector(255 downto 0) := X"E2E1DFDDDBD9D7D6D4D2D0CECCCBC9C7C5C3C2C0BEBCBAB8B7B5B3B1AFADACAA";
constant INIT_H_AVIN_64 : bit_vector(255 downto 0) := X"1717171717171717171717171717171717161616161616161616161616161616";
constant INIT_L_AVIN_64 : bit_vector(255 downto 0) := X"1D1B1918161412100E0D0B090705030200FEFCFAF8F7F5F3F1EFEDECEAE8E6E4";
constant INIT_H_AVIN_65 : bit_vector(255 downto 0) := X"1717171717171717171717171717171717171717171717171717171717171717";
constant INIT_L_AVIN_65 : bit_vector(255 downto 0) := X"58565452504F4D4B4947454442403E3C3A39373533312F2E2C2A28262423211F";
constant INIT_H_AVIN_66 : bit_vector(255 downto 0) := X"1717171717171717171717171717171717171717171717171717171717171717";
constant INIT_L_AVIN_66 : bit_vector(255 downto 0) := X"92908F8D8B8987858482807E7C7A7977757371706E6C6A68666563615F5D5B5A";
constant INIT_H_AVIN_67 : bit_vector(255 downto 0) := X"1717171717171717171717171717171717171717171717171717171717171717";
constant INIT_L_AVIN_67 : bit_vector(255 downto 0) := X"CDCBC9C7C6C4C2C0BEBCBBB9B7B5B3B1B0AEACAAA8A6A5A3A19F9D9B9A989694";
constant INIT_H_AVIN_68 : bit_vector(255 downto 0) := X"1818181818171717171717171717171717171717171717171717171717171717";
constant INIT_L_AVIN_68 : bit_vector(255 downto 0) := X"0806040200FEFDFBF9F7F5F3F2F0EEECEAE8E7E5E3E1DFDDDCDAD8D6D4D2D1CF";
constant INIT_H_AVIN_69 : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_AVIN_69 : bit_vector(255 downto 0) := X"42403E3D3B3937353332302E2C2A28272523211F1D1C1A18161413110F0D0B09";
constant INIT_H_AVIN_6A : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_AVIN_6A : bit_vector(255 downto 0) := X"7D7B7977757472706E6C6A69676563615F5E5C5A58565453514F4D4B49484644";
constant INIT_H_AVIN_6B : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_AVIN_6B : bit_vector(255 downto 0) := X"B7B6B4B2B0AEACABA9A7A5A3A1A09E9C9A98969593918F8D8B8A88868482807F";
constant INIT_H_AVIN_6C : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_AVIN_6C : bit_vector(255 downto 0) := X"F2F0EEECEBE9E7E5E3E1E0DEDCDAD8D6D5D3D1CFCDCBCAC8C6C4C2C0BFBDBBB9";
constant INIT_H_AVIN_6D : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191918181818181818";
constant INIT_L_AVIN_6D : bit_vector(255 downto 0) := X"2D2B2927252322201E1C1A18171513110F0D0C0A0806040201FFFDFBF9F7F6F4";
constant INIT_H_AVIN_6E : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_AVIN_6E : bit_vector(255 downto 0) := X"67656462605E5C5A59575553514F4E4C4A48464443413F3D3B3938363432302E";
constant INIT_H_AVIN_6F : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_AVIN_6F : bit_vector(255 downto 0) := X"A2A09E9C9A99979593918F8E8C8A88868483817F7D7B7978767472706E6D6B69";
constant INIT_H_AVIN_70 : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_AVIN_70 : bit_vector(255 downto 0) := X"DCDBD9D7D5D3D1D0CECCCAC8C6C5C3C1BFBDBBBAB8B6B4B2B0AFADABA9A7A5A4";
constant INIT_H_AVIN_71 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A19191919191919191919191919191919191919";
constant INIT_L_AVIN_71 : bit_vector(255 downto 0) := X"17151311100E0C0A0807050301FFFDFCFAF8F6F4F2F1EFEDEBE9E7E6E4E2E0DE";
constant INIT_H_AVIN_72 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_AVIN_72 : bit_vector(255 downto 0) := X"52504E4C4A48474543413F3D3C3A38363432312F2D2B2927262422201E1C1B19";
constant INIT_H_AVIN_73 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_AVIN_73 : bit_vector(255 downto 0) := X"8C8A89878583817F7E7C7A78767473716F6D6B6968666462605E5D5B59575553";
constant INIT_H_AVIN_74 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_AVIN_74 : bit_vector(255 downto 0) := X"C7C5C3C1BFBEBCBAB8B6B4B3B1AFADABAAA8A6A4A2A09F9D9B9997959492908E";
constant INIT_H_AVIN_75 : bit_vector(255 downto 0) := X"1B1B1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_AVIN_75 : bit_vector(255 downto 0) := X"0100FEFCFAF8F6F5F3F1EFEDEBEAE8E6E4E2E0DFDDDBD9D7D5D4D2D0CECCCAC9";
constant INIT_H_AVIN_76 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_AVIN_76 : bit_vector(255 downto 0) := X"3C3A38373533312F2D2C2A28262422211F1D1B1917161412100E0C0B09070503";
constant INIT_H_AVIN_77 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_AVIN_77 : bit_vector(255 downto 0) := X"777573716F6D6C6A68666462615F5D5B5958565452504E4D4B4947454342403E";
constant INIT_H_AVIN_78 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_AVIN_78 : bit_vector(255 downto 0) := X"B1AFAEACAAA8A6A4A3A19F9D9B9998969492908E8D8B8987858382807E7C7A78";
constant INIT_H_AVIN_79 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_AVIN_79 : bit_vector(255 downto 0) := X"ECEAE8E6E5E3E1DFDDDBDAD8D6D4D2D0CFCDCBC9C7C5C4C2C0BEBCBAB9B7B5B3";
constant INIT_H_AVIN_7A : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_AVIN_7A : bit_vector(255 downto 0) := X"262523211F1D1B1A18161412100F0D0B090705040200FEFCFBF9F7F5F3F1F0EE";
constant INIT_H_AVIN_7B : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_AVIN_7B : bit_vector(255 downto 0) := X"615F5D5C5A58565452514F4D4B4947464442403E3C3B3937353331302E2C2A28";
constant INIT_H_AVIN_7C : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_AVIN_7C : bit_vector(255 downto 0) := X"9C9A98969493918F8D8B8988868482807E7D7B7977757372706E6C6A68676563";
constant INIT_H_AVIN_7D : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_AVIN_7D : bit_vector(255 downto 0) := X"D6D4D3D1CFCDCBC9C8C6C4C2C0BEBDBBB9B7B5B3B2B0AEACAAA8A7A5A3A19F9E";
constant INIT_H_AVIN_7E : bit_vector(255 downto 0) := X"1D1D1D1D1D1D1D1D1D1D1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_AVIN_7E : bit_vector(255 downto 0) := X"110F0D0B0A0806040200FFFDFBF9F7F5F4F2F0EEECEAE9E7E5E3E1DFDEDCDAD8";
constant INIT_H_AVIN_7F : bit_vector(255 downto 0) := X"1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D";
constant INIT_L_AVIN_7F : bit_vector(255 downto 0) := X"4C4A48464442413F3D3B3937363432302E2C2B2927252321201E1C1A18161513";
constant INIT_H_DVIN_00 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_DVIN_00 : bit_vector(255 downto 0) := X"38363533312F2D2B2A28262422201F1D1B1917151412100E0C0A090705030100";
constant INIT_H_DVIN_01 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_DVIN_01 : bit_vector(255 downto 0) := X"73716F6D6C6A68666462615F5D5B5957565452504E4C4B4947454341403E3C3A";
constant INIT_H_DVIN_02 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_DVIN_02 : bit_vector(255 downto 0) := X"ADACAAA8A6A4A3A19F9D9B9998969492908E8D8B8987858382807E7C7A787775";
constant INIT_H_DVIN_03 : bit_vector(255 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000";
constant INIT_L_DVIN_03 : bit_vector(255 downto 0) := X"E8E6E4E3E1DFDDDBD9D8D6D4D2D0CECDCBC9C7C5C3C2C0BEBCBAB8B7B5B3B1AF";
constant INIT_H_DVIN_04 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101000000000000000000000000";
constant INIT_L_DVIN_04 : bit_vector(255 downto 0) := X"23211F1D1B1A18161412100F0D0B090705040200FEFCFAF9F7F5F3F1EFEEECEA";
constant INIT_H_DVIN_05 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_DVIN_05 : bit_vector(255 downto 0) := X"5D5B5A58565452504F4D4B4947464442403E3C3B3937353331302E2C2A282625";
constant INIT_H_DVIN_06 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_DVIN_06 : bit_vector(255 downto 0) := X"98969492918F8D8B8987868482807E7C7B7977757371706E6C6A68666563615F";
constant INIT_H_DVIN_07 : bit_vector(255 downto 0) := X"0101010101010101010101010101010101010101010101010101010101010101";
constant INIT_L_DVIN_07 : bit_vector(255 downto 0) := X"D3D1CFCDCBC9C8C6C4C2C0BEBDBBB9B7B5B3B2B0AEACAAA8A7A5A3A19F9D9C9A";
constant INIT_H_DVIN_08 : bit_vector(255 downto 0) := X"0202020202020202010101010101010101010101010101010101010101010101";
constant INIT_L_DVIN_08 : bit_vector(255 downto 0) := X"0D0B090806040200FEFDFBF9F7F5F4F2F0EEECEAE9E7E5E3E1DFDEDCDAD8D6D4";
constant INIT_H_DVIN_09 : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_DVIN_09 : bit_vector(255 downto 0) := X"48464442403F3D3B3937353432302E2C2A29272523211F1E1C1A18161413110F";
constant INIT_H_DVIN_0A : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_DVIN_0A : bit_vector(255 downto 0) := X"82817F7D7B7977767472706E6C6B6967656361605E5C5A58565553514F4D4B4A";
constant INIT_H_DVIN_0B : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_DVIN_0B : bit_vector(255 downto 0) := X"BDBBB9B7B6B4B2B0AEACABA9A7A5A3A1A09E9C9A98979593918F8D8C8A888684";
constant INIT_H_DVIN_0C : bit_vector(255 downto 0) := X"0202020202020202020202020202020202020202020202020202020202020202";
constant INIT_L_DVIN_0C : bit_vector(255 downto 0) := X"F8F6F4F2F0EEEDEBE9E7E5E3E2E0DEDCDAD8D7D5D3D1CFCDCCCAC8C6C4C2C1BF";
constant INIT_H_DVIN_0D : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030302020202";
constant INIT_L_DVIN_0D : bit_vector(255 downto 0) := X"32302F2D2B2927252422201E1C1A19171513110F0E0C0A0806040301FFFDFBF9";
constant INIT_H_DVIN_0E : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_DVIN_0E : bit_vector(255 downto 0) := X"6D6B6967656462605E5C5A59575553514F4E4C4A48464443413F3D3B3A383634";
constant INIT_H_DVIN_0F : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_DVIN_0F : bit_vector(255 downto 0) := X"A7A6A4A2A09E9C9B9997959391908E8C8A88868583817F7D7B7A78767472706F";
constant INIT_H_DVIN_10 : bit_vector(255 downto 0) := X"0303030303030303030303030303030303030303030303030303030303030303";
constant INIT_L_DVIN_10 : bit_vector(255 downto 0) := X"E2E0DEDDDBD9D7D5D3D2D0CECCCAC8C7C5C3C1BFBDBCBAB8B6B4B2B1AFADABA9";
constant INIT_H_DVIN_11 : bit_vector(255 downto 0) := X"0404040404040404040404040404040403030303030303030303030303030303";
constant INIT_L_DVIN_11 : bit_vector(255 downto 0) := X"1D1B1917151312100E0C0A0807050301FFFDFCFAF8F6F4F2F1EFEDEBE9E8E6E4";
constant INIT_H_DVIN_12 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_DVIN_12 : bit_vector(255 downto 0) := X"57555452504E4C4A49474543413F3E3C3A38363433312F2D2B2928262422201E";
constant INIT_H_DVIN_13 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_DVIN_13 : bit_vector(255 downto 0) := X"92908E8C8B8987858381807E7C7A78767573716F6D6B6A68666462605F5D5B59";
constant INIT_H_DVIN_14 : bit_vector(255 downto 0) := X"0404040404040404040404040404040404040404040404040404040404040404";
constant INIT_L_DVIN_14 : bit_vector(255 downto 0) := X"CCCBC9C7C5C3C1C0BEBCBAB8B6B5B3B1AFADABAAA8A6A4A2A09F9D9B99979594";
constant INIT_H_DVIN_15 : bit_vector(255 downto 0) := X"0505050505040404040404040404040404040404040404040404040404040404";
constant INIT_L_DVIN_15 : bit_vector(255 downto 0) := X"0705030200FEFCFAF8F7F5F3F1EFEDECEAE8E6E4E2E1DFDDDBD9D7D6D4D2D0CE";
constant INIT_H_DVIN_16 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_DVIN_16 : bit_vector(255 downto 0) := X"42403E3C3A38373533312F2E2C2A28262423211F1D1B1918161412100E0D0B09";
constant INIT_H_DVIN_17 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_DVIN_17 : bit_vector(255 downto 0) := X"7C7A79777573716F6E6C6A68666463615F5D5B5958565452504E4D4B49474543";
constant INIT_H_DVIN_18 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_DVIN_18 : bit_vector(255 downto 0) := X"B7B5B3B1B0AEACAAA8A6A5A3A19F9D9B9A98969492908F8D8B8987858482807E";
constant INIT_H_DVIN_19 : bit_vector(255 downto 0) := X"0505050505050505050505050505050505050505050505050505050505050505";
constant INIT_L_DVIN_19 : bit_vector(255 downto 0) := X"F1F0EEECEAE8E6E5E3E1DFDDDCDAD8D6D4D2D1CFCDCBC9C7C6C4C2C0BEBCBBB9";
constant INIT_H_DVIN_1A : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060605050505050505";
constant INIT_L_DVIN_1A : bit_vector(255 downto 0) := X"2C2A28272523211F1D1C1A18161412110F0D0B090706040200FEFCFBF9F7F5F3";
constant INIT_H_DVIN_1B : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_DVIN_1B : bit_vector(255 downto 0) := X"676563615F5E5C5A58565453514F4D4B4948464442403E3D3B3937353332302E";
constant INIT_H_DVIN_1C : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_DVIN_1C : bit_vector(255 downto 0) := X"A19F9E9C9A98969493918F8D8B8988868482807F7D7B7977757472706E6C6A69";
constant INIT_H_DVIN_1D : bit_vector(255 downto 0) := X"0606060606060606060606060606060606060606060606060606060606060606";
constant INIT_L_DVIN_1D : bit_vector(255 downto 0) := X"DCDAD8D6D5D3D1CFCDCBCAC8C6C4C2C0BFBDBBB9B7B5B4B2B0AEACAAA9A7A5A3";
constant INIT_H_DVIN_1E : bit_vector(255 downto 0) := X"0707070707070707070707070706060606060606060606060606060606060606";
constant INIT_L_DVIN_1E : bit_vector(255 downto 0) := X"171513110F0D0C0A0806040201FFFDFBF9F7F6F4F2F0EEECEBE9E7E5E3E1E0DE";
constant INIT_H_DVIN_1F : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_DVIN_1F : bit_vector(255 downto 0) := X"514F4D4C4A48464442413F3D3B3937363432302E2C2B2927252322201E1C1A18";
constant INIT_H_DVIN_20 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_DVIN_20 : bit_vector(255 downto 0) := X"8C8A88868483817F7D7B7978767472706E6D6B6967656362605E5C5A58575553";
constant INIT_H_DVIN_21 : bit_vector(255 downto 0) := X"0707070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_DVIN_21 : bit_vector(255 downto 0) := X"C6C5C3C1BFBDBBBAB8B6B4B2B0AFADABA9A7A5A4A2A09E9C9A99979593918F8E";
constant INIT_H_DVIN_22 : bit_vector(255 downto 0) := X"0807070707070707070707070707070707070707070707070707070707070707";
constant INIT_L_DVIN_22 : bit_vector(255 downto 0) := X"01FFFDFBFAF8F6F4F2F0EFEDEBE9E7E5E4E2E0DEDCDAD9D7D5D3D1D0CECCCAC8";
constant INIT_H_DVIN_23 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_DVIN_23 : bit_vector(255 downto 0) := X"3C3A38363432312F2D2B2927262422201E1C1B1917151311100E0C0A08060503";
constant INIT_H_DVIN_24 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_DVIN_24 : bit_vector(255 downto 0) := X"767473716F6D6B6968666462605E5D5B5957555352504E4C4A48474543413F3D";
constant INIT_H_DVIN_25 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_DVIN_25 : bit_vector(255 downto 0) := X"B1AFADABA9A8A6A4A2A09E9D9B9997959392908E8C8A88878583817F7D7C7A78";
constant INIT_H_DVIN_26 : bit_vector(255 downto 0) := X"0808080808080808080808080808080808080808080808080808080808080808";
constant INIT_L_DVIN_26 : bit_vector(255 downto 0) := X"EBEAE8E6E4E2E0DFDDDBD9D7D5D4D2D0CECCCAC9C7C5C3C1BFBEBCBAB8B6B4B3";
constant INIT_H_DVIN_27 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090908080808080808080808";
constant INIT_L_DVIN_27 : bit_vector(255 downto 0) := X"262422201F1D1B1917161412100E0C0B090705030100FEFCFAF8F6F5F3F1EFED";
constant INIT_H_DVIN_28 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_DVIN_28 : bit_vector(255 downto 0) := X"615F5D5B5957565452504E4C4B4947454341403E3C3A38363533312F2D2B2A28";
constant INIT_H_DVIN_29 : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_DVIN_29 : bit_vector(255 downto 0) := X"9B9998969492908E8D8B8987858382807E7C7A78777573716F6D6C6A68666462";
constant INIT_H_DVIN_2A : bit_vector(255 downto 0) := X"0909090909090909090909090909090909090909090909090909090909090909";
constant INIT_L_DVIN_2A : bit_vector(255 downto 0) := X"D6D4D2D0CECDCBC9C7C5C4C2C0BEBCBAB9B7B5B3B1AFAEACAAA8A6A4A3A19F9D";
constant INIT_H_DVIN_2B : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A09090909090909090909090909090909090909090909";
constant INIT_L_DVIN_2B : bit_vector(255 downto 0) := X"100F0D0B090705040200FEFCFAF9F7F5F3F1EFEEECEAE8E6E4E3E1DFDDDBD9D8";
constant INIT_H_DVIN_2C : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_DVIN_2C : bit_vector(255 downto 0) := X"4B4947464442403E3C3B3937353331302E2C2A28262523211F1D1B1A18161412";
constant INIT_H_DVIN_2D : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_DVIN_2D : bit_vector(255 downto 0) := X"868482807E7C7B7977757371706E6C6A68676563615F5D5C5A58565452514F4D";
constant INIT_H_DVIN_2E : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_DVIN_2E : bit_vector(255 downto 0) := X"C0BEBDBBB9B7B5B3B2B0AEACAAA8A7A5A3A19F9D9C9A98969492918F8D8B8987";
constant INIT_H_DVIN_2F : bit_vector(255 downto 0) := X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A";
constant INIT_L_DVIN_2F : bit_vector(255 downto 0) := X"FBF9F7F5F4F2F0EEECEAE9E7E5E3E1DFDEDCDAD8D6D4D3D1CFCDCBC9C8C6C4C2";
constant INIT_H_DVIN_30 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0A0A";
constant INIT_L_DVIN_30 : bit_vector(255 downto 0) := X"353432302E2C2A29272523211F1E1C1A18161413110F0D0B0A0806040200FFFD";
constant INIT_H_DVIN_31 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_DVIN_31 : bit_vector(255 downto 0) := X"706E6C6B6967656361605E5C5A58565553514F4D4B4A48464442403F3D3B3937";
constant INIT_H_DVIN_32 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_DVIN_32 : bit_vector(255 downto 0) := X"ABA9A7A5A3A2A09E9C9A98979593918F8D8C8A88868482817F7D7B7977767472";
constant INIT_H_DVIN_33 : bit_vector(255 downto 0) := X"0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_DVIN_33 : bit_vector(255 downto 0) := X"E5E3E2E0DEDCDAD8D7D5D3D1CFCDCCCAC8C6C4C2C1BFBDBBB9B8B6B4B2B0AEAD";
constant INIT_H_DVIN_34 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B0B0B0B0B0B0B0B";
constant INIT_L_DVIN_34 : bit_vector(255 downto 0) := X"201E1C1A19171513110F0E0C0A0806040301FFFDFBF9F8F6F4F2F0EEEDEBE9E7";
constant INIT_H_DVIN_35 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_DVIN_35 : bit_vector(255 downto 0) := X"5B5957555351504E4C4A48464543413F3D3B3A38363432302F2D2B2927252422";
constant INIT_H_DVIN_36 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_DVIN_36 : bit_vector(255 downto 0) := X"959391908E8C8A88868583817F7D7B7A78767472706F6D6B6967656462605E5C";
constant INIT_H_DVIN_37 : bit_vector(255 downto 0) := X"0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_DVIN_37 : bit_vector(255 downto 0) := X"D0CECCCAC8C7C5C3C1BFBDBCBAB8B6B4B2B1AFADABA9A7A6A4A2A09E9C9B9997";
constant INIT_H_DVIN_38 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C";
constant INIT_L_DVIN_38 : bit_vector(255 downto 0) := X"0A0807050301FFFEFCFAF8F6F4F3F1EFEDEBE9E8E6E4E2E0DEDDDBD9D7D5D3D2";
constant INIT_H_DVIN_39 : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_DVIN_39 : bit_vector(255 downto 0) := X"4543413F3E3C3A38363433312F2D2B2928262422201E1D1B1917151312100E0C";
constant INIT_H_DVIN_3A : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_DVIN_3A : bit_vector(255 downto 0) := X"807E7C7A78767573716F6D6B6A68666462605F5D5B5957555452504E4C4A4947";
constant INIT_H_DVIN_3B : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_DVIN_3B : bit_vector(255 downto 0) := X"BAB8B6B5B3B1AFADACAAA8A6A4A2A19F9D9B9997969492908E8C8B8987858381";
constant INIT_H_DVIN_3C : bit_vector(255 downto 0) := X"0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D";
constant INIT_L_DVIN_3C : bit_vector(255 downto 0) := X"F5F3F1EFEDECEAE8E6E4E2E1DFDDDBD9D7D6D4D2D0CECCCBC9C7C5C3C1C0BEBC";
constant INIT_H_DVIN_3D : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0D0D0D0D0D";
constant INIT_L_DVIN_3D : bit_vector(255 downto 0) := X"2F2E2C2A28262423211F1D1B1918161412100E0D0B090705030200FEFCFAF8F7";
constant INIT_H_DVIN_3E : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_DVIN_3E : bit_vector(255 downto 0) := X"6A68666463615F5D5B5958565452504F4D4B4947454442403E3C3A3937353331";
constant INIT_H_DVIN_3F : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_DVIN_3F : bit_vector(255 downto 0) := X"A5A3A19F9D9B9A98969492908F8D8B8987858482807E7C7A79777573716F6E6C";
constant INIT_H_DVIN_40 : bit_vector(255 downto 0) := X"0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_DVIN_40 : bit_vector(255 downto 0) := X"DFDDDCDAD8D6D4D2D1CFCDCBC9C7C6C4C2C0BEBCBBB9B7B5B3B1B0AEACAAA8A6";
constant INIT_H_DVIN_41 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E";
constant INIT_L_DVIN_41 : bit_vector(255 downto 0) := X"1A18161412110F0D0B090706040200FEFCFBF9F7F5F3F2F0EEECEAE8E7E5E3E1";
constant INIT_H_DVIN_42 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_DVIN_42 : bit_vector(255 downto 0) := X"5453514F4D4B4948464442403E3D3B3937353332302E2C2A28272523211F1D1C";
constant INIT_H_DVIN_43 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_DVIN_43 : bit_vector(255 downto 0) := X"8F8D8B8A88868482807F7D7B7977757472706E6C6A69676563615F5E5C5A5856";
constant INIT_H_DVIN_44 : bit_vector(255 downto 0) := X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_DVIN_44 : bit_vector(255 downto 0) := X"CAC8C6C4C2C0BFBDBBB9B7B5B4B2B0AEACAAA9A7A5A3A1A09E9C9A9896959391";
constant INIT_H_DVIN_45 : bit_vector(255 downto 0) := X"1010100F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F";
constant INIT_L_DVIN_45 : bit_vector(255 downto 0) := X"040201FFFDFBF9F7F6F4F2F0EEECEBE9E7E5E3E1E0DEDCDAD8D6D5D3D1CFCDCB";
constant INIT_H_DVIN_46 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_DVIN_46 : bit_vector(255 downto 0) := X"3F3D3B3938363432302E2D2B2927252322201E1C1A18171513110F0D0C0A0806";
constant INIT_H_DVIN_47 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_DVIN_47 : bit_vector(255 downto 0) := X"7978767472706E6D6B6967656362605E5C5A58575553514F4D4C4A4846444341";
constant INIT_H_DVIN_48 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_DVIN_48 : bit_vector(255 downto 0) := X"B4B2B0AFADABA9A7A5A4A2A09E9C9A99979593918F8E8C8A88868483817F7D7B";
constant INIT_H_DVIN_49 : bit_vector(255 downto 0) := X"1010101010101010101010101010101010101010101010101010101010101010";
constant INIT_L_DVIN_49 : bit_vector(255 downto 0) := X"EFEDEBE9E7E6E4E2E0DEDCDBD9D7D5D3D1D0CECCCAC8C6C5C3C1BFBDBBBAB8B6";
constant INIT_H_DVIN_4A : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111101010101010101010";
constant INIT_L_DVIN_4A : bit_vector(255 downto 0) := X"2927262422201E1C1B1917151311100E0C0A0806050301FFFDFBFAF8F6F4F2F0";
constant INIT_H_DVIN_4B : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_DVIN_4B : bit_vector(255 downto 0) := X"6462605E5D5B5957555352504E4C4A48474543413F3D3C3A38363432312F2D2B";
constant INIT_H_DVIN_4C : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_DVIN_4C : bit_vector(255 downto 0) := X"9E9D9B9997959492908E8C8A89878583817F7E7C7A78767473716F6D6B696866";
constant INIT_H_DVIN_4D : bit_vector(255 downto 0) := X"1111111111111111111111111111111111111111111111111111111111111111";
constant INIT_L_DVIN_4D : bit_vector(255 downto 0) := X"D9D7D5D4D2D0CECCCAC9C7C5C3C1BFBEBCBAB8B6B4B3B1AFADABA9A8A6A4A2A0";
constant INIT_H_DVIN_4E : bit_vector(255 downto 0) := X"1212121212121212121212121111111111111111111111111111111111111111";
constant INIT_L_DVIN_4E : bit_vector(255 downto 0) := X"1412100E0C0B090705030100FEFCFAF8F6F5F3F1EFEDEBEAE8E6E4E2E0DFDDDB";
constant INIT_H_DVIN_4F : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_DVIN_4F : bit_vector(255 downto 0) := X"4E4C4B4947454341403E3C3A38373533312F2D2C2A28262422211F1D1B191716";
constant INIT_H_DVIN_50 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_DVIN_50 : bit_vector(255 downto 0) := X"8987858382807E7C7A78777573716F6D6C6A68666462615F5D5B595756545250";
constant INIT_H_DVIN_51 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_DVIN_51 : bit_vector(255 downto 0) := X"C4C2C0BEBCBAB9B7B5B3B1AFAEACAAA8A6A4A3A19F9D9B9998969492908E8D8B";
constant INIT_H_DVIN_52 : bit_vector(255 downto 0) := X"1212121212121212121212121212121212121212121212121212121212121212";
constant INIT_L_DVIN_52 : bit_vector(255 downto 0) := X"FEFCFAF9F7F5F3F1EFEEECEAE8E6E4E3E1DFDDDBDAD8D6D4D2D0CFCDCBC9C7C5";
constant INIT_H_DVIN_53 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_DVIN_53 : bit_vector(255 downto 0) := X"3937353331302E2C2A28262523211F1D1B1A18161412100F0D0B090705040200";
constant INIT_H_DVIN_54 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_DVIN_54 : bit_vector(255 downto 0) := X"7372706E6C6A68676563615F5D5C5A58565452514F4D4B4947464442403E3C3B";
constant INIT_H_DVIN_55 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_DVIN_55 : bit_vector(255 downto 0) := X"AEACAAA8A7A5A3A19F9D9C9A98969492918F8D8B8988868482807E7D7B797775";
constant INIT_H_DVIN_56 : bit_vector(255 downto 0) := X"1313131313131313131313131313131313131313131313131313131313131313";
constant INIT_L_DVIN_56 : bit_vector(255 downto 0) := X"E9E7E5E3E1DFDEDCDAD8D6D4D3D1CFCDCBC9C8C6C4C2C0BEBDBBB9B7B5B3B2B0";
constant INIT_H_DVIN_57 : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414131313131313131313131313";
constant INIT_L_DVIN_57 : bit_vector(255 downto 0) := X"2321201E1C1A18161513110F0D0B0A0806040200FFFDFBF9F7F5F4F2F0EEECEA";
constant INIT_H_DVIN_58 : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_DVIN_58 : bit_vector(255 downto 0) := X"5E5C5A58565553514F4D4B4A48464442403F3D3B3937353432302E2C2B292725";
constant INIT_H_DVIN_59 : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_DVIN_59 : bit_vector(255 downto 0) := X"98979593918F8D8C8A88868482817F7D7B7977767472706E6C6B696765636160";
constant INIT_H_DVIN_5A : bit_vector(255 downto 0) := X"1414141414141414141414141414141414141414141414141414141414141414";
constant INIT_L_DVIN_5A : bit_vector(255 downto 0) := X"D3D1CFCECCCAC8C6C4C3C1BFBDBBB9B8B6B4B2B0AEADABA9A7A5A3A2A09E9C9A";
constant INIT_H_DVIN_5B : bit_vector(255 downto 0) := X"1515151515151515141414141414141414141414141414141414141414141414";
constant INIT_L_DVIN_5B : bit_vector(255 downto 0) := X"0E0C0A0806040301FFFDFBF9F8F6F4F2F0EEEDEBE9E7E5E3E2E0DEDCDAD8D7D5";
constant INIT_H_DVIN_5C : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_DVIN_5C : bit_vector(255 downto 0) := X"48464543413F3D3B3A38363432302F2D2B2927252422201E1C1A19171513110F";
constant INIT_H_DVIN_5D : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_DVIN_5D : bit_vector(255 downto 0) := X"83817F7D7C7A78767472716F6D6B6967666462605E5C5B5957555351504E4C4A";
constant INIT_H_DVIN_5E : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_DVIN_5E : bit_vector(255 downto 0) := X"BDBCBAB8B6B4B2B1AFADABA9A7A6A4A2A09E9C9B9997959391908E8C8A888685";
constant INIT_H_DVIN_5F : bit_vector(255 downto 0) := X"1515151515151515151515151515151515151515151515151515151515151515";
constant INIT_L_DVIN_5F : bit_vector(255 downto 0) := X"F8F6F4F3F1EFEDEBE9E8E6E4E2E0DEDDDBD9D7D5D3D2D0CECCCAC8C7C5C3C1BF";
constant INIT_H_DVIN_60 : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161615151515";
constant INIT_L_DVIN_60 : bit_vector(255 downto 0) := X"33312F2D2B2928262422201F1D1B1917151412100E0C0A0907050301FFFEFCFA";
constant INIT_H_DVIN_61 : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161616161616";
constant INIT_L_DVIN_61 : bit_vector(255 downto 0) := X"6D6B6A68666462605F5D5B5957555452504E4C4A49474543413F3E3C3A383634";
constant INIT_H_DVIN_62 : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161616161616";
constant INIT_L_DVIN_62 : bit_vector(255 downto 0) := X"A8A6A4A2A19F9D9B9997969492908E8C8B8987858381807E7C7A78767573716F";
constant INIT_H_DVIN_63 : bit_vector(255 downto 0) := X"1616161616161616161616161616161616161616161616161616161616161616";
constant INIT_L_DVIN_63 : bit_vector(255 downto 0) := X"E2E1DFDDDBD9D7D6D4D2D0CECCCBC9C7C5C3C2C0BEBCBAB8B7B5B3B1AFADACAA";
constant INIT_H_DVIN_64 : bit_vector(255 downto 0) := X"1717171717171717171717171717171717161616161616161616161616161616";
constant INIT_L_DVIN_64 : bit_vector(255 downto 0) := X"1D1B1918161412100E0D0B090705030200FEFCFAF8F7F5F3F1EFEDECEAE8E6E4";
constant INIT_H_DVIN_65 : bit_vector(255 downto 0) := X"1717171717171717171717171717171717171717171717171717171717171717";
constant INIT_L_DVIN_65 : bit_vector(255 downto 0) := X"58565452504F4D4B4947454442403E3C3A39373533312F2E2C2A28262423211F";
constant INIT_H_DVIN_66 : bit_vector(255 downto 0) := X"1717171717171717171717171717171717171717171717171717171717171717";
constant INIT_L_DVIN_66 : bit_vector(255 downto 0) := X"92908F8D8B8987858482807E7C7A7977757371706E6C6A68666563615F5D5B5A";
constant INIT_H_DVIN_67 : bit_vector(255 downto 0) := X"1717171717171717171717171717171717171717171717171717171717171717";
constant INIT_L_DVIN_67 : bit_vector(255 downto 0) := X"CDCBC9C7C6C4C2C0BEBCBBB9B7B5B3B1B0AEACAAA8A6A5A3A19F9D9B9A989694";
constant INIT_H_DVIN_68 : bit_vector(255 downto 0) := X"1818181818171717171717171717171717171717171717171717171717171717";
constant INIT_L_DVIN_68 : bit_vector(255 downto 0) := X"0806040200FEFDFBF9F7F5F3F2F0EEECEAE8E7E5E3E1DFDDDCDAD8D6D4D2D1CF";
constant INIT_H_DVIN_69 : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_DVIN_69 : bit_vector(255 downto 0) := X"42403E3D3B3937353332302E2C2A28272523211F1D1C1A18161413110F0D0B09";
constant INIT_H_DVIN_6A : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_DVIN_6A : bit_vector(255 downto 0) := X"7D7B7977757472706E6C6A69676563615F5E5C5A58565453514F4D4B49484644";
constant INIT_H_DVIN_6B : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_DVIN_6B : bit_vector(255 downto 0) := X"B7B6B4B2B0AEACABA9A7A5A3A1A09E9C9A98969593918F8D8B8A88868482807F";
constant INIT_H_DVIN_6C : bit_vector(255 downto 0) := X"1818181818181818181818181818181818181818181818181818181818181818";
constant INIT_L_DVIN_6C : bit_vector(255 downto 0) := X"F2F0EEECEBE9E7E5E3E1E0DEDCDAD8D6D5D3D1CFCDCBCAC8C6C4C2C0BFBDBBB9";
constant INIT_H_DVIN_6D : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191918181818181818";
constant INIT_L_DVIN_6D : bit_vector(255 downto 0) := X"2D2B2927252322201E1C1A18171513110F0D0C0A0806040201FFFDFBF9F7F6F4";
constant INIT_H_DVIN_6E : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_DVIN_6E : bit_vector(255 downto 0) := X"67656462605E5C5A59575553514F4E4C4A48464443413F3D3B3938363432302E";
constant INIT_H_DVIN_6F : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_DVIN_6F : bit_vector(255 downto 0) := X"A2A09E9C9A99979593918F8E8C8A88868483817F7D7B7978767472706E6D6B69";
constant INIT_H_DVIN_70 : bit_vector(255 downto 0) := X"1919191919191919191919191919191919191919191919191919191919191919";
constant INIT_L_DVIN_70 : bit_vector(255 downto 0) := X"DCDBD9D7D5D3D1D0CECCCAC8C6C5C3C1BFBDBBBAB8B6B4B2B0AFADABA9A7A5A4";
constant INIT_H_DVIN_71 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A19191919191919191919191919191919191919";
constant INIT_L_DVIN_71 : bit_vector(255 downto 0) := X"17151311100E0C0A0807050301FFFDFCFAF8F6F4F2F1EFEDEBE9E7E6E4E2E0DE";
constant INIT_H_DVIN_72 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_DVIN_72 : bit_vector(255 downto 0) := X"52504E4C4A48474543413F3D3C3A38363432312F2D2B2927262422201E1C1B19";
constant INIT_H_DVIN_73 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_DVIN_73 : bit_vector(255 downto 0) := X"8C8A89878583817F7E7C7A78767473716F6D6B6968666462605E5D5B59575553";
constant INIT_H_DVIN_74 : bit_vector(255 downto 0) := X"1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_DVIN_74 : bit_vector(255 downto 0) := X"C7C5C3C1BFBEBCBAB8B6B4B3B1AFADABAAA8A6A4A2A09F9D9B9997959492908E";
constant INIT_H_DVIN_75 : bit_vector(255 downto 0) := X"1B1B1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A";
constant INIT_L_DVIN_75 : bit_vector(255 downto 0) := X"0100FEFCFAF8F6F5F3F1EFEDEBEAE8E6E4E2E0DFDDDBD9D7D5D4D2D0CECCCAC9";
constant INIT_H_DVIN_76 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_DVIN_76 : bit_vector(255 downto 0) := X"3C3A38373533312F2D2C2A28262422211F1D1B1917161412100E0C0B09070503";
constant INIT_H_DVIN_77 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_DVIN_77 : bit_vector(255 downto 0) := X"777573716F6D6C6A68666462615F5D5B5958565452504E4D4B4947454342403E";
constant INIT_H_DVIN_78 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_DVIN_78 : bit_vector(255 downto 0) := X"B1AFAEACAAA8A6A4A3A19F9D9B9998969492908E8D8B8987858382807E7C7A78";
constant INIT_H_DVIN_79 : bit_vector(255 downto 0) := X"1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_DVIN_79 : bit_vector(255 downto 0) := X"ECEAE8E6E5E3E1DFDDDBDAD8D6D4D2D0CFCDCBC9C7C5C4C2C0BEBCBAB9B7B5B3";
constant INIT_H_DVIN_7A : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1B1B1B1B1B1B1B1B1B1B";
constant INIT_L_DVIN_7A : bit_vector(255 downto 0) := X"262523211F1D1B1A18161412100F0D0B090705040200FEFCFBF9F7F5F3F1F0EE";
constant INIT_H_DVIN_7B : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_DVIN_7B : bit_vector(255 downto 0) := X"615F5D5C5A58565452514F4D4B4947464442403E3C3B3937353331302E2C2A28";
constant INIT_H_DVIN_7C : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_DVIN_7C : bit_vector(255 downto 0) := X"9C9A98969493918F8D8B8988868482807E7D7B7977757372706E6C6A68676563";
constant INIT_H_DVIN_7D : bit_vector(255 downto 0) := X"1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_DVIN_7D : bit_vector(255 downto 0) := X"D6D4D3D1CFCDCBC9C8C6C4C2C0BEBDBBB9B7B5B3B2B0AEACAAA8A7A5A3A19F9E";
constant INIT_H_DVIN_7E : bit_vector(255 downto 0) := X"1D1D1D1D1D1D1D1D1D1D1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C";
constant INIT_L_DVIN_7E : bit_vector(255 downto 0) := X"110F0D0B0A0806040200FFFDFBF9F7F5F4F2F0EEECEAE9E7E5E3E1DFDEDCDAD8";
constant INIT_H_DVIN_7F : bit_vector(255 downto 0) := X"1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D";
constant INIT_L_DVIN_7F : bit_vector(255 downto 0) := X"4C4A48464442413F3D3B3937363432302E2C2B2927252321201E1C1A18161513";
end SlowAdcPkg;
