-------------------------------------------------------------------------------
-- File       : AppPkg.vhd
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 2017-04-21
-- Last update: 2018-06-22
-------------------------------------------------------------------------------
-- Description: Application's Package File
-------------------------------------------------------------------------------
-- This file is part of 'EPIX HR Firmware'.
-- It is subject to the license terms in the LICENSE.txt file found in the 
-- top-level directory of this distribution and at: 
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html. 
-- No part of 'EPIX HR Firmware', including this file, 
-- may be copied, modified, propagated, or distributed except according to 
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

use work.StdRtlPkg.all;
use work.AxiLitePkg.all;

package AppPkg is


   constant NUMBER_OF_ASICS_C : natural := 1   
   constant NUMBER_OF_LANES_C : natural := 4;   
   
   constant HR_FD_NUM_AXI_MASTER_SLOTS_C  : natural := 20;
   constant HR_FD_NUM_AXI_SLAVE_SLOTS_C   : natural := 1;
   
   constant PLLREGS_AXI_INDEX_C           : natural := 0;
   constant TRIG_REG_AXI_INDEX_C          : natural := 1;
   constant PRBS0_AXI_INDEX_C             : natural := 2;
   constant PRBS1_AXI_INDEX_C             : natural := 3;
   constant PRBS2_AXI_INDEX_C             : natural := 4;
   constant PRBS3_AXI_INDEX_C             : natural := 5;
   constant AXI_STREAM_MON_INDEX_C        : natural := 6;
   constant DDR_MEM_INDEX_C               : natural := 7;
   constant SACIREGS_AXI_INDEX_C          : natural := 8;
   constant POWER_MODULE_INDEX_C          : natural := 9;
   constant DAC8812_REG_AXI_INDEX_C       : natural := 10;
   constant DACWFMEM_REG_AXI_INDEX_C      : natural := 11;
   constant DAC_MODULE_INDEX_C            : natural := 12;
   constant SCOPE_REG_AXI_INDEX_C         : natural := 13;
   constant ADC_RD_AXI_INDEX_C            : natural := 14;   
   constant ADC_CFG_AXI_INDEX_C           : natural := 15;   
   constant MONADC_REG_AXI_INDEX_C        : natural := 16;
   constant EQUALIZER_REG_AXI_INDEX_C     : natural := 17;
   constant PROG_SUPPLY_REG_AXI_INDEX_C   : natural := 18;
   constant CLK_JIT_CLR_REG_AXI_INDEX_C   : natural := 19;
   
   constant PLLREGS_AXI_BASE_ADDR_C         : slv(31 downto 0) := X"00000000";--0
   constant TRIG_REG_AXI_BASE_ADDR_C        : slv(31 downto 0) := X"01000000";--1
   constant PRBS0_AXI_BASE_ADDR_C           : slv(31 downto 0) := X"02000000";--2
   constant PRBS1_AXI_BASE_ADDR_C           : slv(31 downto 0) := X"02100000";--3
   constant PRBS2_AXI_BASE_ADDR_C           : slv(31 downto 0) := X"02200000";--4
   constant PRBS3_AXI_BASE_ADDR_C           : slv(31 downto 0) := X"02300000";--5
   constant AXI_STREAM_MON_BASE_ADDR_C      : slv(31 downto 0) := X"02400000";--6
   constant DDR_MEM_BASE_ADDR_C             : slv(31 downto 0) := X"03000000";--7
   constant SACIREGS_BASE_ADDR_C            : slv(31 downto 0) := X"04000000";--8
   constant POWER_MODULE_BASE_ADDR_C        : slv(31 downto 0) := X"05000000";--9
   constant DAC8812_AXI_BASE_ADDR_C         : slv(31 downto 0) := X"06000000";--10
   constant DACWFMEM_AXI_BASE_ADDR_C        : slv(31 downto 0) := X"06100000";--11
   constant DAC_MODULE_ADDR_C               : slv(31 downto 0) := X"06200000";--12
   constant SCOPE_REG_AXI_ADDR_C            : slv(31 downto 0) := X"07000000";--13
   constant ADC_RD_AXI_ADDR_C               : slv(31 downto 0) := X"08000000";--14
   constant ADC_CFG_AXI_ADDR_C              : slv(31 downto 0) := X"08100000";--15
   constant MONADC_REG_AXI_ADDR_C           : slv(31 downto 0) := X"08200000";--16
   constant EQUALIZER_REG_AXI_ADDR_C        : slv(31 downto 0) := X"09000000";--17
   constant PROG_SUPPLY_REG_AXI_ADDR_C      : slv(31 downto 0) := X"09100000";--18
   constant CLK_JIT_CLR_REG_AXI_ADDR_C      : slv(31 downto 0) := X"09200000";--19
   
   
   constant HR_FD_AXI_CROSSBAR_MASTERS_CONFIG_C : AxiLiteCrossbarMasterConfigArray(HR_FD_NUM_AXI_MASTER_SLOTS_C-1 downto 0) := (
      PLLREGS_AXI_INDEX_C       => (
         baseAddr             => PLLREGS_AXI_BASE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      TRIG_REG_AXI_INDEX_C      => ( 
         baseAddr             => TRIG_REG_AXI_BASE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      PRBS0_AXI_INDEX_C        => ( 
         baseAddr             => PRBS0_AXI_BASE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      PRBS1_AXI_INDEX_C        => ( 
         baseAddr             => PRBS1_AXI_BASE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      PRBS2_AXI_INDEX_C        => ( 
         baseAddr             => PRBS2_AXI_BASE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      PRBS3_AXI_INDEX_C        => ( 
         baseAddr             => PRBS3_AXI_BASE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      AXI_STREAM_MON_INDEX_C   => ( 
         baseAddr             => AXI_STREAM_MON_BASE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      DDR_MEM_INDEX_C          => ( 
         baseAddr             => DDR_MEM_BASE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),      
      SACIREGS_AXI_INDEX_C     => ( 
         baseAddr             => SACIREGS_BASE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),      
      POWER_MODULE_INDEX_C    => ( 
         baseAddr             => POWER_MODULE_BASE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      DAC8812_REG_AXI_INDEX_C      => ( 
         baseAddr             => DAC8812_AXI_BASE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      DACWFMEM_REG_AXI_INDEX_C      => ( 
         baseAddr             => DACWFMEM_AXI_BASE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      DAC_MODULE_INDEX_C            => ( 
         baseAddr             => DAC_MODULE_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      SCOPE_REG_AXI_INDEX_C         => ( 
         baseAddr             => SCOPE_REG_AXI_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
     ADC_RD_AXI_INDEX_C         => ( 
         baseAddr             => ADC_RD_AXI_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      ADC_CFG_AXI_INDEX_C         => ( 
         baseAddr             => ADC_CFG_AXI_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      MONADC_REG_AXI_INDEX_C        => ( 
         baseAddr             => MONADC_REG_AXI_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      EQUALIZER_REG_AXI_INDEX_C        => ( 
         baseAddr             => EQUALIZER_REG_AXI_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      PROG_SUPPLY_REG_AXI_INDEX_C        => ( 
         baseAddr             => PROG_SUPPLY_REG_AXI_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF"),
      CLK_JIT_CLR_REG_AXI_INDEX_C        => ( 
         baseAddr             => CLK_JIT_CLR_REG_AXI_ADDR_C,
         addrBits             => 20,
         connectivity         => x"FFFF")
   );


   type AppConfigType is record
      AppVersion           : slv(31 downto 0);
   end record;


   constant APP_CONFIG_INIT_C : AppConfigType := (
      AppVersion           => (others => '0')
   );
   
   type HR_FDConfigType is record
      pwrEnableReq         : sl;
   end record;

   constant HR_FD_CONFIG_INIT_C : HR_FDConfigType := (
      pwrEnableReq         => '0'
   );
   

end package AppPkg;

package body AppPkg is

end package body AppPkg;
