-------------------------------------------------------------------------------
-- File       : Hr16bAdcDeserializerUS.vhd
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 2016-05-26
-- Last update: 2019-05-08
-------------------------------------------------------------------------------
-- Description:
-- ADC data deserializer
-- Receives serial ADC Data from an Hr12bAdc SLAC ASIC.
-- Designed specifically for Xilinx Ultrascale series FPGAs
-------------------------------------------------------------------------------
-- This file is part of 'SLAC Firmware Standard Library'.
-- It is subject to the license terms in the LICENSE.txt file found in the 
-- top-level directory of this distribution and at: 
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html. 
-- No part of 'SLAC Firmware Standard Library', including this file, 
-- may be copied, modified, propagated, or distributed except according to 
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library UNISIM;
use UNISIM.vcomponents.all;

use work.StdRtlPkg.all;
use work.AxiLitePkg.all;
use work.AxiStreamPkg.all;
use work.HrAdcPkg.all;

entity Hr16bAdcDeserializer is
   generic (
      TPD_G             : time                 := 1 ns;
      NUM_CHANNELS_G    : natural range 1 to 8 := 8;
      IODELAY_GROUP_G   : string               := "DEFAULT_GROUP";
      IDELAYCTRL_FREQ_G : real                 := 350.0;
      DEFAULT_DELAY_G   : slv(8  downto 0)     := (others => '0');
      FRAME_PATTERN_G   : slv(19 downto 0)     := "11111111110000000000";
      ADC_INVERT_CH_G   : sl                   := '0';
      BIT_REV_G         : sl                   := '0';
      MSB_LSB_G         : sl                   := '1' -- '0' for "MSB_FIRST"
                                                      -- and '1' for "LSB_FIRST"
                                                      );
   port (
      -- Reset for adc deserializer
      adcClkRst : in  sl;                -- global reset
      idelayRst : in  sl;                -- register based reset  
      iserdesRst: in  sl;                -- register based reset 
      -- Serial Data from ADC
      dClk      : in  sl;                       -- Data clock
      dClkDiv4  : in  sl;
      dClkDiv5  : in  sl;
      sDataP    : in  sl;                       -- Frame clock
      sDataN    : in  sl;
      sDataOutP : out sl;                       -- copy of the data
      sDataOutN : out sl;     
      -- Signal to control data gearboxes
      loadDelay       : in sl;
      delay           : in slv(8 downto 0) := "000000000";
      delayValueOut   : out slv(8 downto 0);
      bitSlip         : in slv(2 downto 0) := "000";
      tenbOrder       : in sl := '1';
      gearboxOffset   : in slv(1 downto 0) := "00";
      dataValid       : out sl;
      tenbData        : out Slv10Array(63 downto 0);            
      pixData         : out slv(19 downto 0)     
      );
end Hr16bAdcDeserializer;

-- Define architecture
architecture rtl of Hr16bAdcDeserializer is

  attribute keep : string;
  -------------------------------------------------------------------------------------------------
  -- ADC Readout Clocked Registers
  -------------------------------------------------------------------------------------------------
  type AdcClkDiv4RegType is record
    masterData         : slv(7  downto 0);
    masterData_1       : slv(7  downto 0);
    longDataCounter    : slv(2  downto 0);
    longData           : slv(39 downto 0);
    longData_1         : slv(39 downto 0);
    bitSlip            : slv(2  downto 0);
    masterDataBS       : slv(7  downto 0);
    masterDataBS_1     : slv(7  downto 0);
    longDataStable     : sl;
  end record;

  constant ADC_CLK_DV4_REG_INIT_C : AdcClkDiv4RegType := (
    masterData         => (others => '0'),
    masterData_1       => (others => '0'),
    longDataCounter    => (others => '0'),
    longData           => (others => '0'),
    longData_1         => (others => '0'),
    bitSlip            => (others => '0'),
    masterDataBS       => (others => '0'),
    masterDataBS_1     => (others => '0'),
    longDataStable     => '0'
    );

  type AdcClkDiv5RegType is record
    gearboxCounter      : slv(1 downto 0);
    gearboxSeq          : slv(1 downto 0);
    tenbData            : Slv10Array(63 downto 0);
    masterPixData       : slv(19 downto 0);
    tenbOrder           : sl;
    dataAligned         : sl;
    valid               : sl;
    pixDataGearboxIn    : slv(7 downto 0);
    pixDataGearboxIn_1  : slv(7 downto 0);
    
  end record;

  constant ADC_CLK_DV5_REG_INIT_C : AdcClkDiv5RegType := (
    gearboxCounter      => (others => '0'),
    gearboxSeq          => (others => '0'),
    tenbData            => (others=>(others=>'0')),
    masterPixData       => (others => '0'),
    tenbOrder           => '0',
    dataAligned         => '0',
    valid               => '0',
    pixDataGearboxIn    => (others => '0'),
    pixDataGearboxIn_1  => (others => '0')
    );

  
  
  signal adcDV4R   : AdcClkDiv4RegType := ADC_CLK_DV4_REG_INIT_C;
  signal adcDv4Rin : AdcClkDiv4RegType;

  signal adcDV5R   : AdcClkDiv5RegType := ADC_CLK_DV5_REG_INIT_C;
  signal adcDv5Rin : AdcClkDiv5RegType;
  

   -- Local signals
  signal sDataPadP  : sl;
  signal sDataPadN  : sl;
  signal sData_i    : sl;
  signal sData_d    : sl;

  -- iserdes signal
  signal masterData      : slv(7 downto 0);

  attribute keep of adcDV4R          : signal is "true";
  attribute keep of adcDV5R          : signal is "true";
  attribute keep of sData_i          : signal is "true";

begin

  PixData <= adcDv5R.masterPixData(10)&adcDv5R.masterPixData(11)&adcDv5R.masterPixData(12)&adcDv5R.masterPixData(13)&adcDv5R.masterPixData(14)&adcDv5R.masterPixData(15)&adcDv5R.masterPixData(16)&adcDv5R.masterPixData(17)&adcDv5R.masterPixData(18)&adcDv5R.masterPixData(19)&adcDv5R.masterPixData(0)&adcDv5R.masterPixData(1)&adcDv5R.masterPixData(2)&adcDv5R.masterPixData(3)&adcDv5R.masterPixData(4)&adcDv5R.masterPixData(5)&adcDv5R.masterPixData(6)&adcDv5R.masterPixData(7)&adcDv5R.masterPixData(8)&adcDv5R.masterPixData(9)                       when BIT_REV_G = '1'
             else adcDv5R.masterPixData;

  sDataOutP <= sDataPadP;
  sDataOutN <= sDataPadN;
  -------------------------------------------------------------------------------------------------
  -- Create Clocks
  -------------------------------------------------------------------------------------------------
  
  -- input sData buffer
  --
  U_IBUFDS_sData : IBUFDS_DIFF_OUT
    generic map (
      DQS_BIAS => "FALSE"  -- (FALSE, TRUE)
      )
    port map (
      O  => sDataPadP,   -- 1-bit output: Buffer output
      OB => sDataPadN,
      I  => sDataP,   -- 1-bit input: Diff_p buffer input (connect directly to top-level port)
      IB => sDataN  -- 1-bit input: Diff_n buffer input (connect directly to top-level port)
      );
  -- Optionally invert the pad input
  sData_i <= sDataPadP when ADC_INVERT_CH_G = '0' else sDataPadN;
  ----------------------------------------------------------------------------
  -- idelay3 
  ----------------------------------------------------------------------------
  U_IDELAYE3_0 : IDELAYE3
    generic map (
      CASCADE => "NONE",          -- Cascade setting (MASTER, NONE, SLAVE_END, SLAVE_MIDDLE)
      DELAY_FORMAT => "COUNT",     -- Units of the DELAY_VALUE (COUNT, TIME)
      DELAY_SRC => "IDATAIN",     -- Delay input (DATAIN, IDATAIN)
      DELAY_TYPE => "VAR_LOAD",   -- Set the type of tap delay line (FIXED, VARIABLE, VAR_LOAD)
      DELAY_VALUE => conv_integer(DEFAULT_DELAY_G), -- Input delay value setting
      IS_CLK_INVERTED => '0',     -- Optional inversion for CLK
      IS_RST_INVERTED => '0',     -- Optional inversion for RST
      REFCLK_FREQUENCY => IDELAYCTRL_FREQ_G,  -- IDELAYCTRL clock input frequency in MHz (200.0-2667.0)
      SIM_DEVICE => "ULTRASCALE", -- Set the device version (ULTRASCALE, ULTRASCALE_PLUS, ULTRASCALE_PLUS_ES1,
                                  -- ULTRASCALE_PLUS_ES2)
      UPDATE_MODE => "ASYNC"      -- Determines when updates to the delay will take effect (ASYNC, MANUAL,
                                  -- SYNC)
      )
    port map (
      CASC_OUT => OPEN,       -- 1-bit output: Cascade delay output to ODELAY input cascade
      CNTVALUEOUT => delayValueOut, -- 9-bit output: Counter value output
      DATAOUT => sData_d,         -- 1-bit output: Delayed data output
      CASC_IN => '1',         -- 1-bit input: Cascade delay input from slave ODELAY CASCADE_OUT
      CASC_RETURN => '1', -- 1-bit input: Cascade delay returning from slave ODELAY DATAOUT
      CE => '0',                   -- 1-bit input: Active high enable increment/decrement input
      CLK => dClkDiv4,                 -- 1-bit input: Clock input
      CNTVALUEIN => delay,   -- 9-bit input: Counter value input
      DATAIN => '1',           -- 1-bit input: Data input from the logic
      EN_VTC => '0',           -- 1-bit input: Keep delay constant over VT
      IDATAIN => sData_i,         -- 1-bit input: Data input from the IOBUF
      INC => '0',                 -- 1-bit input: Increment / Decrement tap delay input
      LOAD => loadDelay,               -- 1-bit input: Load DELAY_VALUE input
      RST => idelayRst            -- 1-bit input: Asynchronous Reset to the DELAY_VALUE
      );    
   
  ----------------------------------------------------------------------------
  -- iserdes3
  ----------------------------------------------------------------------------
  U_ISERDESE3_master : ISERDESE3
    generic map (
      DATA_WIDTH => 8,            -- Parallel data width (4,8)
      FIFO_ENABLE => "FALSE",     -- Enables the use of the FIFO
      FIFO_SYNC_MODE => "FALSE",  -- Enables the use of internal 2-stage synchronizers on the FIFO
      IS_CLK_B_INVERTED => '1',   -- Optional inversion for CLK_B
      IS_CLK_INVERTED => '0',     -- Optional inversion for CLK
      IS_RST_INVERTED => '0',     -- Optional inversion for RST
      SIM_DEVICE => "ULTRASCALE"  -- Set the device version (ULTRASCALE, ULTRASCALE_PLUS, ULTRASCALE_PLUS_ES1,
                                  -- ULTRASCALE_PLUS_ES2)
      )
    port map (
      FIFO_EMPTY => OPEN,         -- 1-bit output: FIFO empty flag
      INTERNAL_DIVCLK => open,    -- 1-bit output: Internally divided down clock used when FIFO is
                                  -- disabled (do not connect)

      Q => masterData,            -- bit registered output
      CLK => dClk,            -- 1-bit input: High-speed clock
      CLKDIV => dClkDiv4,         -- 1-bit input: Divided Clock
      CLK_B => dClk,        -- 1-bit input: Inversion of High-speed clock CLK
      D => sData_d,               -- 1-bit input: Serial Data Input
      FIFO_RD_CLK => '1',         -- 1-bit input: FIFO read clock
      FIFO_RD_EN => '1',          -- 1-bit input: Enables reading the FIFO when asserted
      RST => iserdesRst           -- 1-bit input: Asynchronous Reset
      );

  -----------------------------------------------------------------------------
  -- custom logic 
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  -- 8 to 16, 56 gearbox and bitSlip control logic
  -- Part or all 56 bits can be used for idelay3 adjustment
  -----------------------------------------------------------------------------
  adc8to56GearboxComb : process (adcDv4R, masterData, bitSlip) is
    variable v : AdcClkDiv4RegType;
  begin

     v := adcDv4R;

     -- update register with signal values
     v.masterData   := masterData;
     v.bitSlip      := bitSlip;

     -- creates pipeline
     v.masterData_1 := adcDv4R.masterData;
     v.longData_1   := adcDv4R.longData;
     v.masterDataBS_1 := adcDv4R.masterDataBS;
     
     -- data checks on this logic.
     -- 56 bit assembly logic
     case (adcDv4R.longDataCounter) is
       when "000" =>
         v.longData(7 downto 0) := adcDv4R.masterData_1;
         v.longDataCounter := adcDv4R.longDataCounter + 1;
       when "001" =>
         v.longData(15 downto 8) := adcDv4R.masterData_1;
         v.longDataCounter := adcDv4R.longDataCounter + 1;
       when "010" =>
         v.longData(23 downto 16) := adcDv4R.masterData_1;
         v.longDataCounter := adcDv4R.longDataCounter + 1;
       when "011" =>
         v.longData(31 downto 24) := adcDv4R.masterData_1;
         v.longDataCounter := adcDv4R.longDataCounter + 1;            
       when "100" =>
         v.longData(39 downto 32) := adcDv4R.masterData_1;
         v.longDataCounter := (others => '0');
       when others =>
         v.longData  := (others => '0');
         v.longDataCounter := (others => '0');
     end case;

     if adcDv4R.longDataCounter = "000" then
       if adcDv4r.longData = adcDv4r.longData_1 then
         v.longDataStable := '1';
       else
         v.longDataStable := '0';
       end if;
     end if;
   
     --bit slip logic
     case (adcDv4R.bitSlip) is
       when "000" =>
         v.masterDataBS := adcDv4R.masterData(7 downto 0);
       when "001" =>
         v.masterDataBS := adcDv4R.masterData(6 downto 0) & adcDv4R.masterData_1(7);
       when "010" =>
         v.masterDataBS := adcDv4R.masterData(5 downto 0) & adcDv4R.masterData_1(7 downto 6);
       when "011" =>
         v.masterDataBS := adcDv4R.masterData(4 downto 0) & adcDv4R.masterData_1(7 downto 5);
       when "100" =>
         v.masterDataBS := adcDv4R.masterData(3 downto 0) & adcDv4R.masterData_1(7 downto 4);
       when "101" =>
         v.masterDataBS := adcDv4R.masterData(2 downto 0) & adcDv4R.masterData_1(7 downto 3);
       when "110" =>
         v.masterDataBS := adcDv4R.masterData(1 downto 0) & adcDv4R.masterData_1(7 downto 2);
       when "111" =>
         v.masterDataBS := adcDv4R.masterData(0)          & adcDv4R.masterData_1(7 downto  1);
       when others =>
         v.masterDataBS := (others => '0');
     end case;

     adcDv4Rin <= v;
         
     --outputs
     
   end process;

  adclongSeq : process (adcClkRst, dClkDiv4, adcDv4Rin) is 
  begin
    if (adcClkRst = '1') then           
      adcDv4R <= ADC_CLK_DV4_REG_INIT_C;
    elsif (rising_edge(dClkDiv4)) then
      -- latch deserializer data
      adcDv4R <= adcDv4Rin  after TPD_G;
    end if;      
  end process;
   
          
  adc8To7GearboxComb : process (adcDv4R, adcDv5R, gearboxOffset, tenbOrder) is
    variable v : AdcClkDiv5RegType;
  begin

    v := adcDv5R;

    v.tenbOrder           := tenbOrder;
    v.gearboxSeq          := adcDv5R.gearboxCounter + gearboxOffset;
    v.pixDataGearboxIn    := adcDv4R.masterDataBS;
    v.pixDataGearboxIn_1  := adcDv4R.masterDataBS_1;
    
    -- flag that indicates data, or frame signal matches the expected pattern
    if adcDv5R.masterPixData = FRAME_PATTERN_G then
      v.dataAligned := '1';
    else
      v.dataAligned := '0';
    end if;

    if MSB_LSB_G = '1' then             -- LSB
      case (adcDv5R.gearboxSeq) is
        when "00" =>
          v.tenbData(0)   := adcDv5R.pixDataGearboxIn( 1 downto 0) & adcDv5R.pixDataGearboxIn_1( 7 downto 0);
          v.gearboxCounter  := adcDv5R.gearboxCounter + 1;
        when "01" =>
          v.tenbData(0)   := adcDv5R.pixDataGearboxIn( 3 downto 0) & adcDv5R.pixDataGearboxIn_1( 7 downto 2);
          v.gearboxCounter  := adcDv5R.gearboxCounter + 1;
        when "10" =>
          v.tenbData(0)   := adcDv5R.pixDataGearboxIn( 5 downto 0) & adcDv5R.pixDataGearboxIn_1( 7 downto 4);
          v.gearboxCounter  := adcDv5R.gearboxCounter + 1;
        when "11" =>
          v.tenbData(0)   := adcDv5R.pixDataGearboxIn( 7 downto 0) & adcDv5R.pixDataGearboxIn_1( 7 downto 6);
          v.gearboxCounter  := adcDv5R.gearboxCounter + 1;
        when others =>
          v.tenbData(0)   := (others => '0');
          v.gearboxCounter  := (others => '0');
      end case;
    else
      case (adcDv5R.gearboxSeq) is
        when "11" =>
          v.tenbData(0)   := adcDv5R.pixDataGearboxIn( 1 downto 0) & adcDv5R.pixDataGearboxIn_1( 7 downto 0);
          v.gearboxCounter  := adcDv5R.gearboxCounter + 1;
        when "00" =>
          v.tenbData(0)   := adcDv5R.pixDataGearboxIn( 3 downto 0) & adcDv5R.pixDataGearboxIn_1( 7 downto 2);
          v.gearboxCounter  := adcDv5R.gearboxCounter + 1;
        when "01" =>
          v.tenbData(0)   := adcDv5R.pixDataGearboxIn( 5 downto 0) & adcDv5R.pixDataGearboxIn_1( 7 downto 4);
          v.gearboxCounter  := adcDv5R.gearboxCounter + 1;
        when "10" =>
          v.tenbData(0)   := adcDv5R.pixDataGearboxIn( 7 downto 0) & adcDv5R.pixDataGearboxIn_1( 7 downto 6);
          v.gearboxCounter  := adcDv5R.gearboxCounter + 1;
        when others =>
          v.tenbData(0)   := (others => '0');
          v.gearboxCounter  := (others => '0');
      end case;
    end if;

    -- latch whole double word
    v.valid := not adcDv5R.valid;
    if adcDv5R.valid = '1' then
      if adcDv5R.tenbOrder = '0' then
        v.masterPixData  := adcDv5R.tenbData(3) & adcDv5R.tenbData(2);
      else
        v.masterPixData  := adcDv5R.tenbData(2) & adcDv5R.tenbData(3);
      end if;
    end if;
    
    -- 10 bit words pipeline
    for i in 1 to 63 loop
         v.tenbData(i) := adcDv5R.tenbData(i-1);
    end loop;

    adcDv5Rin <= v;
         
    --outputs
    dataValid <= adcDv5R.valid;
    tenbData  <= adcDv5R.tenbData;
    
  end process;
   
   
  adc8To7GearboxSeq : process (adcClkRst, dClkDiv5, adcDv5Rin) is 
  begin
    if (adcClkRst = '1') then
      adcDv5R <= ADC_CLK_DV5_REG_INIT_C;
    elsif (rising_edge(dClkDiv5)) then
      -- latch deserializer data
      adcDv5R <= adcDv5Rin after TPD_G;
    end if;  
  end process;
end rtl;

